* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt nfet a_216_0 a_n84_0 a_94_0 a_30_620
X0 a_94_0 a_30_620 a_n84_0 a_216_0 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
C0 a_94_0 a_n84_0 0.165958f
C1 a_94_0 a_30_620 0.019538f
C2 a_30_620 a_n84_0 0.019538f
C3 a_94_0 a_216_0 0.390769f
C4 a_n84_0 a_216_0 0.122563f
C5 a_30_620 a_216_0 0.245509f
.ends

.subckt pfet$1 a_28_n136 a_n92_0 a_94_0 w_n230_n138 VSUBS
X0 a_94_0 a_28_n136 a_n92_0 w_n230_n138 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
C0 a_28_n136 a_94_0 0.019294f
C1 a_n92_0 a_28_n136 0.019294f
C2 w_n230_n138 a_94_0 0.347768f
C3 a_n92_0 w_n230_n138 0.030103f
C4 a_n92_0 a_94_0 0.158457f
C5 w_n230_n138 a_28_n136 0.143541f
C6 a_94_0 VSUBS 0.020884f
C7 a_n92_0 VSUBS 0.091748f
C8 a_28_n136 VSUBS 0.107314f
C9 w_n230_n138 VSUBS 1.92682f
.ends

.subckt TOP VDD GND Vout Vin Vctrl
Xnfet_0 GND Vout Vin Vctrl nfet
Xnfet_1 GND m1_n72_480 GND Vctrl nfet
Xpfet$1_0 m1_n72_480 Vout Vin VDD GND pfet$1
Xpfet$1_1 Vctrl m1_n72_480 VDD VDD GND pfet$1
X0 VDD Vctrl.t2 m1_n72_480 VDD pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=0 l=0
X1 Vin Vctrl.t0 Vout GND nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=0 l=0
X2 GND.t1 Vctrl.t1 m1_n72_480 GND.t0 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=0 l=0
R0 Vctrl.n0 Vctrl.t0 60.5052
R1 Vctrl Vctrl.t2 56.0454
R2 Vctrl.n0 Vctrl.t1 55.9719
R3 Vctrl Vctrl.n0 0.0999737
R4 GND.n0 GND.t0 747.907
R5 GND.n0 GND.t1 2.1605
R6 GND GND.n0 0.00338991
C0 VDD Vout 0.0175f
C1 VDD Vin 0.03091f
C2 Vctrl m1_n72_480 0.984388f
C3 Vin Vout -0.307332f
C4 VDD Vctrl 0.018047f
C5 VDD m1_n72_480 0.303952f
C6 Vctrl Vout 0.674273f
C7 Vin Vctrl 0.768784f
C8 m1_n72_480 Vout 0.625234f
C9 Vin m1_n72_480 0.681179f
C10 Vctrl GND 1.53662f
C11 Vin GND 0.428795f
C12 Vout GND 0.280843f
C13 m1_n72_480 GND 0.441193f
C14 VDD GND 4.089155f
.ends

