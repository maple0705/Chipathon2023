* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt CAP_ARRAY top_c0 top_c1 top_c5 top_c3 top_c2 top_c4 top_c_dummy common_bottom
X0 top_c5.t0 common_bottom.t41 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1 top_c3.t0 common_bottom.t62 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2 top_c5.t1 common_bottom.t40 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3 top_c3.t1 common_bottom.t5 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4 top_c4.t0 common_bottom.t58 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X5 top_c5.t2 common_bottom.t39 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X6 top_c5.t3 common_bottom.t38 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X7 top_c5.t4 common_bottom.t37 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X8 top_c5.t5 common_bottom.t36 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X9 top_c1.t0 common_bottom.t59 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X10 top_c5.t6 common_bottom.t35 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X11 top_c3.t2 common_bottom.t46 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X12 top_c5.t7 common_bottom.t34 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X13 top_c3.t3 common_bottom.t1 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X14 top_c5.t8 common_bottom.t33 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X15 top_c5.t9 common_bottom.t32 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X16 top_c2.t0 common_bottom.t63 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X17 top_c5.t10 common_bottom.t31 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X18 top_c4.t1 common_bottom.t52 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X19 top_c3.t4 common_bottom.t42 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X20 top_c4.t2 common_bottom.t51 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X21 top_c5.t11 common_bottom.t30 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X22 top_c5.t12 common_bottom.t29 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X23 top_c5.t13 common_bottom.t28 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X24 top_c4.t3 common_bottom.t50 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X25 top_c4.t4 common_bottom.t9 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X26 top_c4.t5 common_bottom.t4 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X27 top_c5.t14 common_bottom.t27 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X28 top_c5.t15 common_bottom.t26 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X29 top_c4.t6 common_bottom.t45 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X30 top_c4.t7 common_bottom.t49 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X31 top_c5.t16 common_bottom.t25 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X32 top_c5.t17 common_bottom.t24 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X33 top_c5.t18 common_bottom.t23 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X34 top_c4.t8 common_bottom.t8 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X35 top_c2.t1 common_bottom.t55 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X36 top_c4.t9 common_bottom.t3 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X37 top_c5.t19 common_bottom.t22 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X38 top_c_dummy.t0 common_bottom.t60 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X39 top_c5.t20 common_bottom.t21 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X40 top_c2.t2 common_bottom.t54 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X41 top_c5.t21 common_bottom.t20 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X42 top_c1.t1 common_bottom.t56 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X43 top_c5.t22 common_bottom.t19 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X44 top_c4.t10 common_bottom.t44 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X45 top_c5.t23 common_bottom.t18 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X46 top_c0.t0 common_bottom.t61 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X47 top_c5.t24 common_bottom.t17 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X48 top_c4.t11 common_bottom.t57 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X49 top_c4.t12 common_bottom.t48 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X50 top_c5.t25 common_bottom.t16 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X51 top_c3.t5 common_bottom.t47 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X52 top_c4.t13 common_bottom.t7 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X53 top_c4.t14 common_bottom.t2 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X54 top_c5.t26 common_bottom.t15 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X55 top_c5.t27 common_bottom.t14 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X56 top_c3.t6 common_bottom.t6 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X57 top_c4.t15 common_bottom.t43 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X58 top_c5.t28 common_bottom.t13 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X59 top_c5.t29 common_bottom.t12 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X60 top_c5.t30 common_bottom.t11 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X61 top_c3.t7 common_bottom.t0 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X62 top_c2.t3 common_bottom.t53 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X63 top_c5.t31 common_bottom.t10 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
R0 top_c5.n59 top_c5.n58 47.7474
R1 top_c5.n26 top_c5.n9 10.9803
R2 top_c5.n58 top_c5.n47 6.64175
R3 top_c5.n47 top_c5.n46 5.8095
R4 top_c5.n58 top_c5.n57 4.33906
R5 top_c5.n47 top_c5.n29 4.31121
R6 top_c5.n26 top_c5.n25 4.31121
R7 top_c5.n27 top_c5.n1 4.31121
R8 top_c5.n28 top_c5.n0 4.31121
R9 top_c5.n27 top_c5.n26 3.26675
R10 top_c5.n28 top_c5.n27 3.26675
R11 top_c5.n59 top_c5.n28 2.51225
R12 top_c5.n6 top_c5.n5 1.13669
R13 top_c5.n51 top_c5.n49 0.988357
R14 top_c5.n49 top_c5.n48 0.988357
R15 top_c5.n36 top_c5.n35 0.988357
R16 top_c5.n38 top_c5.n35 0.988357
R17 top_c5.n41 top_c5.n34 0.988357
R18 top_c5.n43 top_c5.n34 0.988357
R19 top_c5.n33 top_c5.n31 0.988357
R20 top_c5.n12 top_c5.n11 0.988357
R21 top_c5.n14 top_c5.n11 0.988357
R22 top_c5.n17 top_c5.n10 0.988357
R23 top_c5.n19 top_c5.n10 0.988357
R24 top_c5.n24 top_c5.n23 0.988357
R25 top_c5.n3 top_c5.n2 0.988357
R26 top_c5.n5 top_c5.n3 0.988357
R27 top_c5.n8 top_c5.n2 0.9777
R28 top_c5.n56 top_c5.n48 0.9605
R29 top_c5.n54 top_c5.n51 0.9605
R30 top_c5.n30 top_c5.n29 0.9605
R31 top_c5.n44 top_c5.n33 0.9605
R32 top_c5.n1 top_c5.n0 0.9605
R33 top_c5.n23 top_c5.n21 0.9605
R34 top_c5.n25 top_c5.n1 0.9605
R35 top_c5.n6 top_c5.t18 0.892022
R36 top_c5.n36 top_c5.t2 0.72448
R37 top_c5.n12 top_c5.t5 0.72448
R38 top_c5.n40 top_c5.n39 0.6605
R39 top_c5.n16 top_c5.n15 0.6605
R40 top_c5.n53 top_c5.n52 0.646689
R41 top_c5.n54 top_c5.n53 0.632643
R42 top_c5.n57 top_c5.n56 0.632643
R43 top_c5.n39 top_c5.n38 0.632643
R44 top_c5.n41 top_c5.n40 0.632643
R45 top_c5.n15 top_c5.n14 0.632643
R46 top_c5.n17 top_c5.n16 0.632643
R47 top_c5.n9 top_c5.n8 0.631
R48 top_c5.n44 top_c5.n43 0.604786
R49 top_c5.n21 top_c5.n19 0.604786
R50 top_c5.n46 top_c5.n45 0.595021
R51 top_c5.n52 top_c5.t25 0.586765
R52 top_c5 top_c5.n59 0.494375
R53 top_c5.n46 top_c5.n30 0.323104
R54 top_c5.n7 top_c5.n6 0.203778
R55 top_c5.n52 top_c5.t10 0.106765
R56 top_c5.n53 top_c5.t23 0.0923367
R57 top_c5.n49 top_c5.t11 0.0923367
R58 top_c5.n50 top_c5.t26 0.0923367
R59 top_c5.n55 top_c5.t12 0.0923367
R60 top_c5.n57 top_c5.t29 0.0923367
R61 top_c5.n35 top_c5.t8 0.0923367
R62 top_c5.n37 top_c5.t24 0.0923367
R63 top_c5.n39 top_c5.t13 0.0923367
R64 top_c5.n40 top_c5.t27 0.0923367
R65 top_c5.n34 top_c5.t28 0.0923367
R66 top_c5.n42 top_c5.t14 0.0923367
R67 top_c5.n31 top_c5.t30 0.0923367
R68 top_c5.n32 top_c5.t16 0.0923367
R69 top_c5.n45 top_c5.t0 0.0923367
R70 top_c5.n11 top_c5.t7 0.0923367
R71 top_c5.n13 top_c5.t22 0.0923367
R72 top_c5.n15 top_c5.t1 0.0923367
R73 top_c5.n16 top_c5.t15 0.0923367
R74 top_c5.n10 top_c5.t31 0.0923367
R75 top_c5.n18 top_c5.t17 0.0923367
R76 top_c5.n20 top_c5.t4 0.0923367
R77 top_c5.n22 top_c5.t20 0.0923367
R78 top_c5.n24 top_c5.t6 0.0923367
R79 top_c5.n3 top_c5.t21 0.0923367
R80 top_c5.n4 top_c5.t3 0.0923367
R81 top_c5.n7 top_c5.t19 0.0923367
R82 top_c5.n9 top_c5.t9 0.0923367
R83 top_c5.n50 top_c5.n48 0.0283571
R84 top_c5.n51 top_c5.n50 0.0283571
R85 top_c5.n56 top_c5.n55 0.0283571
R86 top_c5.n55 top_c5.n54 0.0283571
R87 top_c5.n38 top_c5.n37 0.0283571
R88 top_c5.n37 top_c5.n36 0.0283571
R89 top_c5.n43 top_c5.n42 0.0283571
R90 top_c5.n42 top_c5.n41 0.0283571
R91 top_c5.n31 top_c5.n29 0.0283571
R92 top_c5.n32 top_c5.n30 0.0283571
R93 top_c5.n33 top_c5.n32 0.0283571
R94 top_c5.n45 top_c5.n44 0.0283571
R95 top_c5.n13 top_c5.n12 0.0283571
R96 top_c5.n14 top_c5.n13 0.0283571
R97 top_c5.n18 top_c5.n17 0.0283571
R98 top_c5.n19 top_c5.n18 0.0283571
R99 top_c5.n21 top_c5.n20 0.0283571
R100 top_c5.n20 top_c5.n0 0.0283571
R101 top_c5.n23 top_c5.n22 0.0283571
R102 top_c5.n22 top_c5.n1 0.0283571
R103 top_c5.n25 top_c5.n24 0.0283571
R104 top_c5.n5 top_c5.n4 0.0283571
R105 top_c5.n4 top_c5.n2 0.0283571
R106 top_c5.n8 top_c5.n7 0.0162308
R107 common_bottom common_bottom.t9 6.59189
R108 common_bottom.t7 common_bottom.t1 1.23983
R109 common_bottom.t1 common_bottom.t39 1.23983
R110 common_bottom.t39 common_bottom.t17 1.23983
R111 common_bottom.t17 common_bottom.t28 1.23983
R112 common_bottom.t14 common_bottom.t28 1.23983
R113 common_bottom.t27 common_bottom.t14 1.23983
R114 common_bottom.t47 common_bottom.t36 1.23216
R115 common_bottom.t54 common_bottom.t30 1.23216
R116 common_bottom.t15 common_bottom.t46 1.23216
R117 common_bottom.t29 common_bottom.t18 1.23216
R118 common_bottom.t6 common_bottom.t63 1.23216
R119 common_bottom.t50 common_bottom.t48 1.23216
R120 common_bottom.t42 common_bottom.t13 1.23216
R121 common_bottom.t36 common_bottom.t19 1.23216
R122 common_bottom.t19 common_bottom.t40 1.23216
R123 common_bottom.t34 common_bottom.t3 1.23216
R124 common_bottom.t61 common_bottom.t58 1.23216
R125 common_bottom.t31 common_bottom.t60 1.23216
R126 common_bottom.t16 common_bottom.t59 1.23216
R127 common_bottom.t2 common_bottom.t33 1.23216
R128 common_bottom.t33 common_bottom.t55 1.23216
R129 common_bottom.t26 common_bottom.t24 1.23216
R130 common_bottom.t24 common_bottom.t37 1.23216
R131 common_bottom.t21 common_bottom.t10 1.23216
R132 common_bottom.t35 common_bottom.t8 1.23216
R133 common_bottom.t44 common_bottom.t5 1.23216
R134 common_bottom.t32 common_bottom.t22 1.23216
R135 common_bottom.t57 common_bottom.t38 1.23216
R136 common_bottom.t52 common_bottom.t20 1.23216
R137 common_bottom.t41 common_bottom.t27 1.23216
R138 common_bottom.t47 common_bottom.t30 1.2245
R139 common_bottom.t15 common_bottom.t30 1.2245
R140 common_bottom.t15 common_bottom.t29 1.2245
R141 common_bottom.t29 common_bottom.t6 1.2245
R142 common_bottom.t6 common_bottom.t50 1.2245
R143 common_bottom.t13 common_bottom.t50 1.2245
R144 common_bottom.t13 common_bottom.t27 1.2245
R145 common_bottom.t3 common_bottom.t40 1.2245
R146 common_bottom.t58 common_bottom.t3 1.2245
R147 common_bottom.t60 common_bottom.t58 1.2245
R148 common_bottom.t59 common_bottom.t60 1.2245
R149 common_bottom.t56 common_bottom.t59 1.2245
R150 common_bottom.t42 common_bottom.t14 1.2245
R151 common_bottom.t42 common_bottom.t48 1.2245
R152 common_bottom.t48 common_bottom.t63 1.2245
R153 common_bottom.t63 common_bottom.t18 1.2245
R154 common_bottom.t18 common_bottom.t46 1.2245
R155 common_bottom.t46 common_bottom.t54 1.2245
R156 common_bottom.t36 common_bottom.t54 1.2245
R157 common_bottom.t19 common_bottom.t34 1.2245
R158 common_bottom.t34 common_bottom.t54 1.2245
R159 common_bottom.t34 common_bottom.t61 1.2245
R160 common_bottom.t61 common_bottom.t46 1.2245
R161 common_bottom.t61 common_bottom.t31 1.2245
R162 common_bottom.t31 common_bottom.t18 1.2245
R163 common_bottom.t31 common_bottom.t16 1.2245
R164 common_bottom.t16 common_bottom.t63 1.2245
R165 common_bottom.t51 common_bottom.t56 1.2245
R166 common_bottom.t16 common_bottom.t51 1.2245
R167 common_bottom.t51 common_bottom.t48 1.2245
R168 common_bottom.t2 common_bottom.t28 1.2245
R169 common_bottom.t51 common_bottom.t2 1.2245
R170 common_bottom.t2 common_bottom.t42 1.2245
R171 common_bottom.t33 common_bottom.t17 1.2245
R172 common_bottom.t33 common_bottom.t56 1.2245
R173 common_bottom.t55 common_bottom.t39 1.2245
R174 common_bottom.t55 common_bottom.t62 1.2245
R175 common_bottom.t62 common_bottom.t56 1.2245
R176 common_bottom.t62 common_bottom.t23 1.2245
R177 common_bottom.t23 common_bottom.t59 1.2245
R178 common_bottom.t23 common_bottom.t53 1.2245
R179 common_bottom.t53 common_bottom.t5 1.2245
R180 common_bottom.t53 common_bottom.t60 1.2245
R181 common_bottom.t53 common_bottom.t49 1.2245
R182 common_bottom.t49 common_bottom.t58 1.2245
R183 common_bottom.t49 common_bottom.t0 1.2245
R184 common_bottom.t0 common_bottom.t3 1.2245
R185 common_bottom.t0 common_bottom.t26 1.2245
R186 common_bottom.t26 common_bottom.t40 1.2245
R187 common_bottom.t37 common_bottom.t21 1.2245
R188 common_bottom.t24 common_bottom.t10 1.2245
R189 common_bottom.t0 common_bottom.t10 1.2245
R190 common_bottom.t8 common_bottom.t5 1.2245
R191 common_bottom.t10 common_bottom.t8 1.2245
R192 common_bottom.t49 common_bottom.t8 1.2245
R193 common_bottom.t21 common_bottom.t35 1.2245
R194 common_bottom.t35 common_bottom.t44 1.2245
R195 common_bottom.t32 common_bottom.t57 1.2245
R196 common_bottom.t44 common_bottom.t32 1.2245
R197 common_bottom.t5 common_bottom.t22 1.2245
R198 common_bottom.t23 common_bottom.t22 1.2245
R199 common_bottom.t22 common_bottom.t38 1.2245
R200 common_bottom.t62 common_bottom.t38 1.2245
R201 common_bottom.t1 common_bottom.t20 1.2245
R202 common_bottom.t38 common_bottom.t20 1.2245
R203 common_bottom.t55 common_bottom.t20 1.2245
R204 common_bottom.t57 common_bottom.t52 1.2245
R205 common_bottom.t52 common_bottom.t7 1.2245
R206 common_bottom.t25 common_bottom.t41 1.2245
R207 common_bottom.t13 common_bottom.t25 1.2245
R208 common_bottom.t25 common_bottom.t11 1.2245
R209 common_bottom.t11 common_bottom.t50 1.2245
R210 common_bottom.t11 common_bottom.t45 1.2245
R211 common_bottom.t45 common_bottom.t6 1.2245
R212 common_bottom.t45 common_bottom.t12 1.2245
R213 common_bottom.t12 common_bottom.t29 1.2245
R214 common_bottom.t12 common_bottom.t4 1.2245
R215 common_bottom.t4 common_bottom.t15 1.2245
R216 common_bottom.t4 common_bottom.t43 1.2245
R217 common_bottom.t30 common_bottom.t43 1.2245
R218 common_bottom.t9 common_bottom.t43 1.2245
R219 common_bottom.t9 common_bottom.t47 1.2245
R220 top_c3.n6 top_c3.n5 24.4219
R221 top_c3.n3 top_c3.t4 11.1293
R222 top_c3.n0 top_c3.t3 11.1224
R223 top_c3.n1 top_c3.n0 6.64613
R224 top_c3.n2 top_c3.n1 6.64484
R225 top_c3.n4 top_c3.n3 6.64282
R226 top_c3.n5 top_c3.n4 6.64282
R227 top_c3.n6 top_c3.n2 5.28119
R228 top_c3.n0 top_c3.t0 4.67797
R229 top_c3.n2 top_c3.t7 4.67599
R230 top_c3.n3 top_c3.t6 4.67077
R231 top_c3.n5 top_c3.t5 4.67077
R232 top_c3.n4 top_c3.t2 4.48695
R233 top_c3.n1 top_c3.t1 4.47901
R234 top_c3 top_c3.n6 1.0805
R235 top_c4.n30 top_c4.n29 30.758
R236 top_c4.n29 top_c4.n28 9.81496
R237 top_c4.n22 top_c4.n21 9.81479
R238 top_c4.n23 top_c4.n16 9.7865
R239 top_c4.n24 top_c4.n15 9.7865
R240 top_c4.n26 top_c4.n14 9.7865
R241 top_c4.n27 top_c4.n13 9.7865
R242 top_c4.n7 top_c4.n6 9.44428
R243 top_c4.n4 top_c4.n1 9.416
R244 top_c4.n5 top_c4.n0 9.416
R245 top_c4.n30 top_c4.n12 8.94864
R246 top_c4.n20 top_c4.n19 7.66414
R247 top_c4.n21 top_c4.n20 5.95628
R248 top_c4.n8 top_c4.n7 5.94959
R249 top_c4.n2 top_c4.n1 5.36384
R250 top_c4.n20 top_c4.t6 4.65484
R251 top_c4.n12 top_c4.n11 4.57893
R252 top_c4.n8 top_c4.t10 4.47101
R253 top_c4.n12 top_c4.n8 3.26797
R254 top_c4.n16 top_c4.n15 1.8905
R255 top_c4.n14 top_c4.n13 1.8905
R256 top_c4.n1 top_c4.n0 1.8905
R257 top_c4.n21 top_c4.n16 1.4855
R258 top_c4.n15 top_c4.n14 1.4855
R259 top_c4.n29 top_c4.n13 1.4855
R260 top_c4.n7 top_c4.n0 1.4855
R261 top_c4 top_c4.n30 0.8105
R262 top_c4.n19 top_c4.n18 0.6605
R263 top_c4.n11 top_c4.n10 0.6605
R264 top_c4.n18 top_c4.n17 0.646689
R265 top_c4.n10 top_c4.n9 0.646689
R266 top_c4.n17 top_c4.t14 0.586765
R267 top_c4.n9 top_c4.t9 0.586765
R268 top_c4.n27 top_c4.n26 0.483929
R269 top_c4.n24 top_c4.n23 0.483929
R270 top_c4.n5 top_c4.n4 0.483929
R271 top_c4.n2 top_c4.t13 0.313204
R272 top_c4.n3 top_c4.n2 0.306937
R273 top_c4.n17 top_c4.t2 0.106765
R274 top_c4.n9 top_c4.t0 0.106765
R275 top_c4.n28 top_c4.t4 0.0964127
R276 top_c4.n25 top_c4.t15 0.0923367
R277 top_c4.n22 top_c4.t5 0.0923367
R278 top_c4.n18 top_c4.t12 0.0923367
R279 top_c4.n19 top_c4.t3 0.0923367
R280 top_c4.n10 top_c4.t7 0.0923367
R281 top_c4.n11 top_c4.t8 0.0923367
R282 top_c4.n6 top_c4.t11 0.0923367
R283 top_c4.n3 top_c4.t1 0.0923367
R284 top_c4.n28 top_c4.n27 0.0289832
R285 top_c4.n25 top_c4.n24 0.0287857
R286 top_c4.n26 top_c4.n25 0.0287857
R287 top_c4.n23 top_c4.n22 0.0287857
R288 top_c4.n6 top_c4.n5 0.0287857
R289 top_c4.n4 top_c4.n3 0.0287857
R290 top_c1 top_c1.n0 16.4063
R291 top_c1.n0 top_c1.t1 7.74631
R292 top_c1.n0 top_c1.t0 4.47901
R293 top_c2.n2 top_c2.n1 21.2881
R294 top_c2.n1 top_c2.t0 14.5021
R295 top_c2.n0 top_c2.t1 14.4963
R296 top_c2.n2 top_c2.n0 11.7141
R297 top_c2.n1 top_c2.t2 4.48671
R298 top_c2.n0 top_c2.t3 4.47901
R299 top_c2 top_c2.n2 1.37413
R300 top_c_dummy top_c_dummy.t0 17.575
R301 top_c0 top_c0.t0 14.1362
C0 m3_16090_37400 top_c5 0.577918f
C1 top_c2 top_c5 2.08451f
C2 common_bottom m3_13080_37400 1.11323f
C3 top_c1 top_c5 0.827905f
C4 top_c2 top_c1 0.089709f
C5 top_c_dummy top_c5 0.58041f
C6 common_bottom m3_n1905_37400 0.979483f
C7 top_c2 top_c_dummy 3.45141f
C8 top_c1 top_c_dummy 0.545203f
C9 common_bottom m3_9610_37600 0.974327f
C10 top_c4 m3_13080_37400 0.17303f
C11 common_bottom top_c4 17.2234f
C12 top_c3 m3_13080_37400 3.56255f
C13 top_c3 common_bottom 10.2294f
C14 common_bottom m3_1090_37400 0.975713f
C15 common_bottom top_c0 2.01468f
C16 top_c4 m3_n1905_37400 3.33282f
C17 top_c3 m3_n1905_37400 0.24292f
C18 top_c4 m3_9610_37600 0.283401f
C19 top_c3 m3_9610_37600 0.026205f
C20 top_c3 top_c4 4.8107f
C21 m3_9610_37600 top_c0 0.132431f
C22 m3_13080_37400 top_c5 0.787868f
C23 m3_16090_37400 common_bottom 0.97451f
C24 common_bottom top_c5 31.515802f
C25 top_c4 m3_1090_37400 0.148711f
C26 top_c4 top_c0 0.425447f
C27 top_c2 m3_13080_37400 0.029803f
C28 top_c2 common_bottom 6.59935f
C29 top_c3 m3_1090_37400 3.37214f
C30 top_c3 top_c0 0.171906f
C31 common_bottom top_c1 3.06981f
C32 top_c5 m3_n1905_37400 0.707599f
C33 common_bottom top_c_dummy 1.99712f
C34 m3_9610_37600 top_c5 0.664815f
C35 m3_16090_37400 top_c4 3.72826f
C36 top_c2 m3_9610_37600 3.18787f
C37 top_c4 top_c5 8.70553f
C38 top_c3 m3_16090_37400 0.01917f
C39 top_c2 top_c4 0.731677f
C40 top_c3 top_c5 2.85677f
C41 top_c2 top_c3 2.92517f
C42 m3_1090_37400 top_c5 0.423352f
C43 top_c0 top_c5 1.02447f
C44 top_c2 m3_1090_37400 0.26486f
C45 top_c2 top_c0 0.0776f
C46 top_c4 top_c1 0.426536f
C47 top_c3 top_c1 0.171911f
C48 top_c1 top_c0 3.29281f
C49 top_c4 top_c_dummy 0.484191f
C50 top_c3 top_c_dummy 0.083598f
C51 top_c_dummy top_c0 0.013195f
C52 common_bottom VSUBS 81.923294f
C53 top_c0 VSUBS 7.462662f
C54 top_c1 VSUBS 9.781748f
C55 top_c_dummy VSUBS 7.799115f
C56 top_c2 VSUBS 19.267962f
C57 top_c3 VSUBS 28.25109f
C58 top_c4 VSUBS 45.17333f
C59 top_c5 VSUBS 85.864395f
C60 m3_16090_37400 VSUBS 4.75247f $ **FLOATING
C61 m3_13080_37400 VSUBS 4.85576f $ **FLOATING
C62 m3_9610_37600 VSUBS 4.70657f $ **FLOATING
C63 m3_1090_37400 VSUBS 4.78423f $ **FLOATING
C64 m3_n1905_37400 VSUBS 4.76133f $ **FLOATING
C65 top_c0.t0 VSUBS 5.10498f
C66 top_c_dummy.t0 VSUBS 2.95832f
C67 top_c2.t1 VSUBS 4.23123f
C68 top_c2.t3 VSUBS 3.72597f
C69 top_c2.n0 VSUBS 1.08459f
C70 top_c2.t0 VSUBS 3.6147f
C71 top_c2.t2 VSUBS 3.72912f
C72 top_c2.n1 VSUBS 0.96196f
C73 top_c2.n2 VSUBS 0.89487f
C74 top_c1.t1 VSUBS 2.69345f
C75 top_c1.t0 VSUBS 2.48754f
C76 top_c1.n0 VSUBS 0.805015f
C77 top_c4.n0 VSUBS 0.067791f
C78 top_c4.n1 VSUBS 0.167882f
C79 top_c4.t13 VSUBS 1.9142f
C80 top_c4.n2 VSUBS 0.457151f
C81 top_c4.t1 VSUBS 1.06757f
C82 top_c4.n3 VSUBS 0.872765f
C83 top_c4.n4 VSUBS 0.396233f
C84 top_c4.n5 VSUBS 0.396233f
C85 top_c4.t11 VSUBS 1.06757f
C86 top_c4.n6 VSUBS 0.733244f
C87 top_c4.n7 VSUBS 0.149347f
C88 top_c4.t10 VSUBS 2.01099f
C89 top_c4.n8 VSUBS 0.207098f
C90 top_c4.t0 VSUBS 1.16577f
C91 top_c4.t9 VSUBS 1.86402f
C92 top_c4.n9 VSUBS 1.1434f
C93 top_c4.t7 VSUBS 1.06757f
C94 top_c4.n10 VSUBS 1.04616f
C95 top_c4.t8 VSUBS 1.06757f
C96 top_c4.n11 VSUBS 1.07261f
C97 top_c4.n12 VSUBS 0.248575f
C98 top_c4.n13 VSUBS 0.069219f
C99 top_c4.n14 VSUBS 0.069219f
C100 top_c4.n15 VSUBS 0.069219f
C101 top_c4.n16 VSUBS 0.069219f
C102 top_c4.t2 VSUBS 1.16577f
C103 top_c4.t14 VSUBS 1.86402f
C104 top_c4.n17 VSUBS 1.1434f
C105 top_c4.t12 VSUBS 1.06757f
C106 top_c4.n18 VSUBS 1.04616f
C107 top_c4.t3 VSUBS 1.06757f
C108 top_c4.n19 VSUBS 1.18806f
C109 top_c4.t6 VSUBS 2.05111f
C110 top_c4.n20 VSUBS 0.417766f
C111 top_c4.n21 VSUBS 0.150996f
C112 top_c4.t5 VSUBS 1.06757f
C113 top_c4.n22 VSUBS 0.75331f
C114 top_c4.n23 VSUBS 0.416331f
C115 top_c4.n24 VSUBS 0.416331f
C116 top_c4.t15 VSUBS 1.06757f
C117 top_c4.n25 VSUBS 0.503285f
C118 top_c4.n26 VSUBS 0.416331f
C119 top_c4.n27 VSUBS 0.448328f
C120 top_c4.t4 VSUBS 1.03165f
C121 top_c4.n28 VSUBS 0.835367f
C122 top_c4.n29 VSUBS 0.496705f
C123 top_c4.n30 VSUBS 0.606739f
C124 top_c3.t3 VSUBS 3.21137f
C125 top_c3.t0 VSUBS 2.97684f
C126 top_c3.n0 VSUBS 0.546008f
C127 top_c3.t1 VSUBS 2.88953f
C128 top_c3.n1 VSUBS 0.428324f
C129 top_c3.t7 VSUBS 2.97636f
C130 top_c3.n2 VSUBS 0.389511f
C131 top_c3.t4 VSUBS 2.96484f
C132 top_c3.t6 VSUBS 3.02964f
C133 top_c3.n3 VSUBS 0.467116f
C134 top_c3.t2 VSUBS 2.91497f
C135 top_c3.n4 VSUBS 0.429217f
C136 top_c3.t5 VSUBS 3.14427f
C137 top_c3.n5 VSUBS 0.773749f
C138 top_c3.n6 VSUBS 0.623065f
C139 common_bottom.t43 VSUBS 1.06159f
C140 common_bottom.t30 VSUBS 1.13747f
C141 common_bottom.t54 VSUBS 1.14036f
C142 common_bottom.t40 VSUBS 1.06015f
C143 common_bottom.t3 VSUBS 1.13747f
C144 common_bottom.t58 VSUBS 1.13747f
C145 common_bottom.t46 VSUBS 1.14036f
C146 common_bottom.t60 VSUBS 1.13747f
C147 common_bottom.t18 VSUBS 1.14036f
C148 common_bottom.t59 VSUBS 1.13747f
C149 common_bottom.t63 VSUBS 1.14036f
C150 common_bottom.t56 VSUBS 1.13891f
C151 common_bottom.t48 VSUBS 1.14036f
C152 common_bottom.t28 VSUBS 1.06159f
C153 common_bottom.t14 VSUBS 1.06159f
C154 common_bottom.t50 VSUBS 1.13747f
C155 common_bottom.t27 VSUBS 1.06015f
C156 common_bottom.t41 VSUBS 0.985713f
C157 common_bottom.t6 VSUBS 1.13747f
C158 common_bottom.t29 VSUBS 1.13747f
C159 common_bottom.t15 VSUBS 1.13747f
C160 common_bottom.t4 VSUBS 1.06159f
C161 common_bottom.t12 VSUBS 1.06159f
C162 common_bottom.t45 VSUBS 1.06159f
C163 common_bottom.t11 VSUBS 1.06159f
C164 common_bottom.t25 VSUBS 1.06159f
C165 common_bottom.t13 VSUBS 1.13747f
C166 common_bottom.t42 VSUBS 1.14036f
C167 common_bottom.t17 VSUBS 1.06159f
C168 common_bottom.t39 VSUBS 1.06159f
C169 common_bottom.t20 VSUBS 1.13747f
C170 common_bottom.t38 VSUBS 1.14036f
C171 common_bottom.t22 VSUBS 1.14036f
C172 common_bottom.t5 VSUBS 1.13747f
C173 common_bottom.t8 VSUBS 1.13747f
C174 common_bottom.t10 VSUBS 1.14036f
C175 common_bottom.t1 VSUBS 1.06159f
C176 common_bottom.t7 VSUBS 0.984269f
C177 common_bottom.t52 VSUBS 1.06304f
C178 common_bottom.t57 VSUBS 1.06015f
C179 common_bottom.t32 VSUBS 1.06015f
C180 common_bottom.t44 VSUBS 1.06304f
C181 common_bottom.t35 VSUBS 1.06304f
C182 common_bottom.t21 VSUBS 1.06015f
C183 common_bottom.t37 VSUBS 0.982824f
C184 common_bottom.t24 VSUBS 1.06448f
C185 common_bottom.t26 VSUBS 1.06015f
C186 common_bottom.t0 VSUBS 1.13891f
C187 common_bottom.t49 VSUBS 1.13891f
C188 common_bottom.t53 VSUBS 1.13891f
C189 common_bottom.t23 VSUBS 1.13891f
C190 common_bottom.t62 VSUBS 1.13891f
C191 common_bottom.t55 VSUBS 1.14036f
C192 common_bottom.t33 VSUBS 1.13891f
C193 common_bottom.t2 VSUBS 1.13747f
C194 common_bottom.t51 VSUBS 1.13891f
C195 common_bottom.t16 VSUBS 1.14036f
C196 common_bottom.t31 VSUBS 1.14036f
C197 common_bottom.t61 VSUBS 1.14036f
C198 common_bottom.t34 VSUBS 1.14036f
C199 common_bottom.t19 VSUBS 1.06448f
C200 common_bottom.t36 VSUBS 1.06159f
C201 common_bottom.t47 VSUBS 1.06015f
C202 common_bottom.t9 VSUBS 1.05373f
C203 top_c5.n0 VSUBS 0.229409f
C204 top_c5.n1 VSUBS 0.256356f
C205 top_c5.n2 VSUBS 0.206256f
C206 top_c5.t18 VSUBS 1.24308f
C207 top_c5.t21 VSUBS 0.660201f
C208 top_c5.n3 VSUBS 0.586645f
C209 top_c5.t3 VSUBS 0.660201f
C210 top_c5.n4 VSUBS 0.306522f
C211 top_c5.n5 VSUBS 0.230247f
C212 top_c5.n6 VSUBS 0.131095f
C213 top_c5.t19 VSUBS 0.660201f
C214 top_c5.n7 VSUBS 0.525227f
C215 top_c5.n8 VSUBS 0.215097f
C216 top_c5.t9 VSUBS 0.660201f
C217 top_c5.n9 VSUBS 0.836149f
C218 top_c5.t31 VSUBS 0.660201f
C219 top_c5.n10 VSUBS 0.59314f
C220 top_c5.t7 VSUBS 0.660201f
C221 top_c5.n11 VSUBS 0.580046f
C222 top_c5.t5 VSUBS 1.21077f
C223 top_c5.n12 VSUBS 0.339481f
C224 top_c5.t22 VSUBS 0.660201f
C225 top_c5.n13 VSUBS 0.306522f
C226 top_c5.n14 VSUBS 0.259494f
C227 top_c5.t1 VSUBS 0.660201f
C228 top_c5.n15 VSUBS 0.689303f
C229 top_c5.t15 VSUBS 0.660201f
C230 top_c5.n16 VSUBS 0.689303f
C231 top_c5.n17 VSUBS 0.260148f
C232 top_c5.t17 VSUBS 0.660201f
C233 top_c5.n18 VSUBS 0.306522f
C234 top_c5.n19 VSUBS 0.250597f
C235 top_c5.t4 VSUBS 0.660201f
C236 top_c5.n20 VSUBS 0.306522f
C237 top_c5.n21 VSUBS 0.246902f
C238 top_c5.t20 VSUBS 0.660201f
C239 top_c5.n22 VSUBS 0.306522f
C240 top_c5.n23 VSUBS 0.186741f
C241 top_c5.t6 VSUBS 0.660201f
C242 top_c5.n24 VSUBS 0.462008f
C243 top_c5.n25 VSUBS 0.205157f
C244 top_c5.n26 VSUBS 0.260607f
C245 top_c5.n27 VSUBS 0.083512f
C246 top_c5.n28 VSUBS 0.071498f
C247 top_c5.n29 VSUBS 0.205157f
C248 top_c5.n30 VSUBS 0.256356f
C249 top_c5.t30 VSUBS 0.660201f
C250 top_c5.n31 VSUBS 0.443284f
C251 top_c5.t16 VSUBS 0.660201f
C252 top_c5.n32 VSUBS 0.306522f
C253 top_c5.n33 VSUBS 0.195898f
C254 top_c5.t28 VSUBS 0.660201f
C255 top_c5.n34 VSUBS 0.580046f
C256 top_c5.t8 VSUBS 0.660201f
C257 top_c5.n35 VSUBS 0.580046f
C258 top_c5.t2 VSUBS 1.26677f
C259 top_c5.n36 VSUBS 0.347616f
C260 top_c5.t24 VSUBS 0.660201f
C261 top_c5.n37 VSUBS 0.306522f
C262 top_c5.n38 VSUBS 0.259494f
C263 top_c5.t13 VSUBS 0.660201f
C264 top_c5.n39 VSUBS 0.689303f
C265 top_c5.t27 VSUBS 0.660201f
C266 top_c5.n40 VSUBS 0.689303f
C267 top_c5.n41 VSUBS 0.259494f
C268 top_c5.t14 VSUBS 0.660201f
C269 top_c5.n42 VSUBS 0.306522f
C270 top_c5.n43 VSUBS 0.25087f
C271 top_c5.n44 VSUBS 0.246902f
C272 top_c5.t0 VSUBS 0.660201f
C273 top_c5.n45 VSUBS 0.550638f
C274 top_c5.n46 VSUBS 0.078776f
C275 top_c5.n47 VSUBS 0.175917f
C276 top_c5.n48 VSUBS 0.219726f
C277 top_c5.t11 VSUBS 0.660201f
C278 top_c5.n49 VSUBS 0.602567f
C279 top_c5.t26 VSUBS 0.660201f
C280 top_c5.n50 VSUBS 0.306522f
C281 top_c5.n51 VSUBS 0.195898f
C282 top_c5.t10 VSUBS 0.720928f
C283 top_c5.t25 VSUBS 1.15273f
C284 top_c5.n52 VSUBS 0.707092f
C285 top_c5.t23 VSUBS 0.660201f
C286 top_c5.n53 VSUBS 0.639402f
C287 top_c5.n54 VSUBS 0.230205f
C288 top_c5.t12 VSUBS 0.660201f
C289 top_c5.n55 VSUBS 0.306522f
C290 top_c5.n56 VSUBS 0.230205f
C291 top_c5.t29 VSUBS 0.660201f
C292 top_c5.n57 VSUBS 0.623386f
C293 top_c5.n58 VSUBS 0.579789f
C294 top_c5.n59 VSUBS 0.476295f
.ends

