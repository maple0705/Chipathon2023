** sch_path: /home/nkimura/sw.sch
.subckt TOP Vctrl VDD Vout Vin GND
*.PININFO Vctrl:I Vin:I Vout:O VDD:I GND:I
M1 Vin net1 Vout VDD pfet_03v3 L=0.28u W=2.8u nf=1 m=1
M2 Vin Vctrl Vout GND nfet_03v3 L=0.28u W=2.8u nf=1 m=1
M3 net1 Vctrl VDD VDD pfet_03v3 L=0.28u W=2.8u nf=1 m=1
M4 net1 Vctrl GND GND nfet_03v3 L=0.28u W=2.8u nf=1 m=1
.ends
 * Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__addf_1 A B CI CO S VDD VNW VPW VSS
M_M51 VSS net9 S VPW nfet_05v0 W=7.1e-07 L=6e-07
M_M46 net9 CI net47 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M45 net42 CI VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M34 CO net7 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M33 VDD net9 S VNW pfet_05v0 W=1.215e-06 L=5e-07
M_M28 net9 CI net29 VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M24 net9 net7 net3 VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M25 net3 A VDD VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M26 VDD B net3 VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M27 net3 CI VDD VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M21 net7 CI net1 VNW pfet_05v0 W=7e-07 L=5e-07
M_M20 net19 B net7 VNW pfet_05v0 W=7e-07 L=5e-07
M_M18 VDD A net19 VNW pfet_05v0 W=7e-07 L=5e-07
M_M17 CO net7 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_M48 net47 B net49 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M41 net9 net7 net42 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M43 net42 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M44 VSS B net42 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M38 net7 CI net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M37 net36 B net7 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M35 VSS A net36 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M30 net29 B net31 VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M23 VDD B net1 VNW pfet_05v0 W=7e-07 L=5e-07
M_M22 net1 A VDD VNW pfet_05v0 W=7e-07 L=5e-07
M_M50 net49 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M40 VSS B net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M39 net5 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M32 net31 A VDD VNW pfet_05v0 W=6.6e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__addf_2 A B CI CO S VDD VNW VPW VSS
M_M51_17 VSS net9 S VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M51 VSS net9 S VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M46 net9 CI net47 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M45 net42 CI VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M34 CO net7 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M34_25 CO net7 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M33_12 VDD net9 S VNW pfet_05v0 W=1.12e-06 L=5e-07
M_M33 VDD net9 S VNW pfet_05v0 W=1.12e-06 L=5e-07
M_M28 net9 CI net29 VNW pfet_05v0 W=6.8e-07 L=5e-07
M_M24 net9 net7 net3 VNW pfet_05v0 W=6.8e-07 L=5e-07
M_M25 net3 A VDD VNW pfet_05v0 W=6.8e-07 L=5e-07
M_M26 VDD B net3 VNW pfet_05v0 W=6.8e-07 L=5e-07
M_M27 net3 CI VDD VNW pfet_05v0 W=6.8e-07 L=5e-07
M_M21 net7 CI net1 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M20 net19 B net7 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M18 VDD A net19 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M17 CO net7 VDD VNW pfet_05v0 W=1.195e-06 L=5e-07
M_M17_23 CO net7 VDD VNW pfet_05v0 W=1.195e-06 L=5e-07
M_M48 net47 B net49 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M41 net9 net7 net42 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M43 net42 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M44 VSS B net42 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M38 net7 CI net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M37 net36 B net7 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M35 VSS A net36 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M30 net29 B net31 VNW pfet_05v0 W=6.8e-07 L=5e-07
M_M23 VDD B net1 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M22 net1 A VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M50 net49 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M40 VSS B net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M39 net5 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M32 net31 A VDD VNW pfet_05v0 W=6.8e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__addf_4 A B CI CO S VDD VNW VPW VSS
M_M51_17_0 VSS net9 S VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M51_18 VSS net9 S VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M51_17 VSS net9 S VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M51 VSS net9 S VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M46 net9 CI net47 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M45 net42 CI VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M34 CO net7 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M34_25 CO net7 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M34_53 CO net7 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M34_25_56 CO net7 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_M33_12_23 VDD net9 S VNW pfet_05v0 W=1.095e-06 L=5e-07
M_M33_34 VDD net9 S VNW pfet_05v0 W=1.095e-06 L=5e-07
M_M33_12 VDD net9 S VNW pfet_05v0 W=1.095e-06 L=5e-07
M_M33 VDD net9 S VNW pfet_05v0 W=1.095e-06 L=5e-07
M_M28 net9 CI net29 VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M24 net9 net7 net3 VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M25 net3 A VDD VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M26 VDD B net3 VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M27 net3 CI VDD VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M21 net7 CI net1 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M20 net19 B net7 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M18 VDD A net19 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M17 CO net7 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_M17_23 CO net7 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_M17_66 CO net7 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_M17_23_46 CO net7 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_M48 net47 B net49 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M41 net9 net7 net42 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M43 net42 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M44 VSS B net42 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M38 net7 CI net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M37 net36 B net7 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M35 VSS A net36 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M30 net29 B net31 VNW pfet_05v0 W=6.6e-07 L=5e-07
M_M23 VDD B net1 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M22 net1 A VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_M50 net49 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M40 VSS B net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M39 net5 A VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_M32 net31 A VDD VNW pfet_05v0 W=6.6e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__addh_1 A B CO S VDD VNW VPW VSS
M_i_2 VSS NCO CO VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_5 net_0 A VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_4 NCO B net_0 VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0 S NS VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_3 VDD NCO CO VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7 NCO A VDD VNW pfet_05v0 W=6.35e-07 L=5e-07
M_i_6 VDD B NCO VNW pfet_05v0 W=6.35e-07 L=5e-07
M_i_11 NS A net_2 VNW pfet_05v0 W=6.35e-07 L=5e-07
M_i_13 VDD NCO NS VNW pfet_05v0 W=6.35e-07 L=5e-07
M_i_1 S NS VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9 NS B net_1 VPW nfet_05v0 W=4.2e-07 L=6e-07
M_i_8 net_1 A NS VPW nfet_05v0 W=4.2e-07 L=6e-07
M_i_10 VSS NCO net_1 VPW nfet_05v0 W=4.2e-07 L=6e-07
M_i_12 net_2 B VDD VNW pfet_05v0 W=6.35e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__addh_2 A B CO S VDD VNW VPW VSS
M_i_2_1 CO NCO VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_2_0 VSS NCO CO VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_5 net_0 A VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_4 NCO B net_0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0_1 S NS VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0_0 VSS NS S VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_3_1 CO NCO VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_3_0 VDD NCO CO VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7 NCO A VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6 VDD B NCO VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_11 NS A net_2 VNW pfet_05v0 W=9.75e-07 L=5e-07
M_i_13 VDD NCO NS VNW pfet_05v0 W=9.75e-07 L=5e-07
M_i_1_1 S NS VDD VNW pfet_05v0 W=9.75e-07 L=5e-07
M_i_1_0 VDD NS S VNW pfet_05v0 W=9.75e-07 L=5e-07
M_i_9 NS B net_1 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_8 net_1 A NS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_10 VSS NCO net_1 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_12 net_2 B VDD VNW pfet_05v0 W=9.75e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__addh_4 A B CO S VDD VNW VPW VSS
M_i_5_1 net_0_0 A VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_1 NCO B net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 net_0_1 B NCO VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_0 VSS A net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10_0 net_1 NCO VSS VPW nfet_05v0 W=6.1e-07 L=6e-07
M_i_8_0 NS A net_1 VPW nfet_05v0 W=6.1e-07 L=6e-07
M_i_9_0 net_1 B NS VPW nfet_05v0 W=6.1e-07 L=6e-07
M_i_9_1 NS B net_1 VPW nfet_05v0 W=6.1e-07 L=6e-07
M_i_8_1 net_1 A NS VPW nfet_05v0 W=6.1e-07 L=6e-07
M_i_10_1 VSS NCO net_1 VPW nfet_05v0 W=6.1e-07 L=6e-07
M_i_2_3 CO NCO VSS VPW nfet_05v0 W=1.05e-06 L=6e-07
M_i_2_2 VSS NCO CO VPW nfet_05v0 W=1.05e-06 L=6e-07
M_i_2_1 CO NCO VSS VPW nfet_05v0 W=1.05e-06 L=6e-07
M_i_2_0 VSS NCO CO VPW nfet_05v0 W=1.05e-06 L=6e-07
M_i_0_3 S NS VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 VSS NS S VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 S NS VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 VSS NS S VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7_1 NCO A VDD VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_6_1 VDD B NCO VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_6_0 NCO B VDD VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_7_0 VDD A NCO VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_13_0 NS NCO VDD VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_11_0 net_2_0 A NS VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_12_0 VDD B net_2_0 VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_12_1 net_2_1 B VDD VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_11_1 NS A net_2_1 VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_13_1 VDD NCO NS VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_3_3 CO NCO VDD VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_3_2 VDD NCO CO VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_3_1 CO NCO VDD VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_3_0 VDD NCO CO VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_1_3 S NS VDD VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_1_2 VDD NS S VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_1_1 S NS VDD VNW pfet_05v0 W=9.9e-07 L=5e-07
M_i_1_0 VDD NS S VNW pfet_05v0 W=9.9e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3 VSS A2 net_0 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_4 Z_neg A1 VDD VNW pfet_05v0 W=6e-07 L=5e-07
M_i_5 VDD A2 Z_neg VNW pfet_05v0 W=6e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_3 VSS A2 net_0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_4 Z_neg A1 VDD VNW pfet_05v0 W=1.07e-06 L=5e-07
M_i_5 VDD A2 Z_neg VNW pfet_05v0 W=1.07e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
M_i_3_1 net_0_1 A2 VSS VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_2_1 Z_neg A1 net_0_1 VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_2_0 net_0_0 A1 Z_neg VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_3_0 VSS A2 net_0_0 VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_0_3 Z Z_neg VSS VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_0_2 VSS Z_neg Z VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_0_1 Z Z_neg VSS VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_0_0 VSS Z_neg Z VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_5_1 Z_neg A2 VDD VNW pfet_05v0 W=1.125e-06 L=5e-07
M_i_4_1 VDD A1 Z_neg VNW pfet_05v0 W=1.125e-06 L=5e-07
M_i_4_0 Z_neg A1 VDD VNW pfet_05v0 W=1.125e-06 L=5e-07
M_i_5_0 VDD A2 Z_neg VNW pfet_05v0 W=1.125e-06 L=5e-07
M_i_1_3 Z Z_neg VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_1_2 VDD Z_neg Z VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_1_1 Z Z_neg VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_1_0 VDD Z_neg Z VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_3 net_1 A2 net_0 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_4 VSS A3 net_1 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_5 VDD A1 Z_neg VNW pfet_05v0 W=5.35e-07 L=5e-07
M_i_6 Z_neg A2 VDD VNW pfet_05v0 W=5.35e-07 L=5e-07
M_i_7 VDD A3 Z_neg VNW pfet_05v0 W=5.35e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_3 net_1 A2 net_0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_4 VSS A3 net_1 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_5 VDD A1 Z_neg VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_6 Z_neg A2 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_7 VDD A3 Z_neg VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
M_i_4_0 net_1_1 A3 VSS VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_3_1 net_0_1 A2 net_1_1 VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_2_1 Z_neg A1 net_0_1 VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_2_0 net_0_0 A1 Z_neg VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_3_0 net_1_0 A2 net_0_0 VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_4_1 VSS A3 net_1_0 VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_0_3 Z Z_neg VSS VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_0_2 VSS Z_neg Z VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_0_1 Z Z_neg VSS VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_0_0 VSS Z_neg Z VPW nfet_05v0 W=7.6e-07 L=6e-07
M_i_7_0 Z_neg A3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_1 VDD A2 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_1 Z_neg A1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_0 VDD A1 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0 Z_neg A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 VDD A3 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=4.2e-07 L=6e-07
M_i_3 net_1 A2 net_0 VPW nfet_05v0 W=4.2e-07 L=6e-07
M_i_4 net_2 A3 net_1 VPW nfet_05v0 W=4.2e-07 L=6e-07
M_i_5 VSS A4 net_2 VPW nfet_05v0 W=4.2e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_6 Z_neg A1 VDD VNW pfet_05v0 W=6e-07 L=5e-07
M_i_7 VDD A2 Z_neg VNW pfet_05v0 W=6e-07 L=5e-07
M_i_8 Z_neg A3 VDD VNW pfet_05v0 W=6e-07 L=5e-07
M_i_9 VDD A4 Z_neg VNW pfet_05v0 W=6e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 net_1 A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4 net_2 A3 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5 VSS A4 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6 Z_neg A1 VDD VNW pfet_05v0 W=8.55e-07 L=5e-07
M_i_7 VDD A2 Z_neg VNW pfet_05v0 W=8.55e-07 L=5e-07
M_i_8 Z_neg A3 VDD VNW pfet_05v0 W=8.55e-07 L=5e-07
M_i_9 VDD A4 Z_neg VNW pfet_05v0 W=8.55e-07 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
M_i_5_1 net_2_1 A4 VSS VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_4_1 net_1_1 A3 net_2_1 VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_3_1 net_0_1 A2 net_1_1 VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_2_1 Z_neg A1 net_0_1 VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_2_0 net_0_0 A1 Z_neg VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_3_0 net_1_0 A2 net_0_0 VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_4_0 net_2_0 A3 net_1_0 VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_5_0 VSS A4 net_2_0 VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_0_3 Z Z_neg VSS VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_0_2 VSS Z_neg Z VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_0_1 Z Z_neg VSS VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_0_0 VSS Z_neg Z VPW nfet_05v0 W=6.45e-07 L=6e-07
M_i_9_1 Z_neg A4 VDD VNW pfet_05v0 W=1.11e-06 L=5e-07
M_i_8_1 VDD A3 Z_neg VNW pfet_05v0 W=1.11e-06 L=5e-07
M_i_7_1 Z_neg A2 VDD VNW pfet_05v0 W=1.11e-06 L=5e-07
M_i_6_1 VDD A1 Z_neg VNW pfet_05v0 W=1.11e-06 L=5e-07
M_i_6_0 Z_neg A1 VDD VNW pfet_05v0 W=1.11e-06 L=5e-07
M_i_7_0 VDD A2 Z_neg VNW pfet_05v0 W=1.11e-06 L=5e-07
M_i_8_0 Z_neg A3 VDD VNW pfet_05v0 W=1.11e-06 L=5e-07
M_i_9_0 VDD A4 Z_neg VNW pfet_05v0 W=1.11e-06 L=5e-07
M_i_1_3 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
D0 VPW I diode_nd2ps_06v0 A=0.2052p P=1.86u
* D1 I VNW diode_pd2nw_06v0 A=0.2052p P=1.86u
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
M_i_1 net_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 VSS B ZN VPW nfet_05v0 W=5.1e-07 L=6e-07
M_i_4 ZN A2 net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_3 net_1 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5 VDD B net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
M_i_2_0 ZN B VSS VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_2_1 VSS B ZN VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_1_0 net_0_0 A2 VSS VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_0_1 ZN A1 net_0_0 VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_0_0 net_0_1 A1 ZN VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_1_1 VSS A2 net_0_1 VPW nfet_05v0 W=7.75e-07 L=6e-07
M_i_5_0 VDD B net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_1 net_1 B VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4_0 ZN A2 net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_3_1 net_1 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_3_0 ZN A1 net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4_1 net_1 A2 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
M_i_1_3 net_0_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 ZN A1 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 net_0_1 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 VSS A2 net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0_2 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0_3 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 VSS A2 net_0_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 ZN B VSS VPW nfet_05v0 W=5.1e-07 L=6e-07
M_i_2_2 VSS B ZN VPW nfet_05v0 W=5.1e-07 L=6e-07
M_i_2_1 ZN B VSS VPW nfet_05v0 W=5.1e-07 L=6e-07
M_i_2_0 VSS B ZN VPW nfet_05v0 W=5.1e-07 L=6e-07
M_i_4_3 ZN A2 net_1 VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_3_3 net_1 A1 ZN VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_3_2 ZN A1 net_1 VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_4_2 net_1 A2 ZN VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_4_1 ZN A2 net_1 VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_3_1 net_1 A1 ZN VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_3_0 ZN A1 net_1 VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_4_0 net_1 A2 ZN VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_5_3 VDD B net_1 VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_5_2 net_1 B VDD VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_5_1 VDD B net_1 VNW pfet_05v0 W=1.2e-06 L=5e-07
M_i_5_0 net_1 B VDD VNW pfet_05v0 W=1.2e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
M_i_3 net_1 B2 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_2 ZN B1 net_1 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0 net_0 A1 ZN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_7 VDD B2 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6 net_2 B1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4 ZN A1 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5 net_2 A2 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
M_i_3_1 net_1_0 B2 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_2_1 ZN B1 net_1_0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_2_0 net_1_1 B1 ZN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_3_0 VSS B2 net_1_1 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_1_1 net_0_0 A2 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0_1 ZN A1 net_0_0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0_0 net_0_1 A1 ZN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_1_0 VSS A2 net_0_1 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_7_1 VDD B2 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_1 net_2 B1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_0 VDD B1 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7_0 net_2 B2 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_1 ZN A2 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4_1 net_2 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4_0 ZN A1 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_0 net_2 A2 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
M_i_3_3 net_1_0 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 ZN B1 net_1_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_1_1 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 VSS B2 net_1_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_1_2 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 ZN B1 net_1_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_1_3 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS B2 net_1_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0_1 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 VSS A2 net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_0_2 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN A1 net_0_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 net_0_3 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 VSS A2 net_0_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7_3 VDD B2 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_3 net_2 B1 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_2 VDD B1 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_2 net_2 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 VDD B2 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 net_2 B1 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 VDD B1 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 net_2 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 ZN A2 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 net_2 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_1 ZN A1 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 net_2 A2 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_2 ZN A2 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_2 net_2 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_3 ZN A1 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_3 net_2 A2 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
M_i_1 net_0 A2 VSS VPW nfet_05v0 W=7.1e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=7.1e-07 L=6e-07
M_i_2 VSS B ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_3 ZN C VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_5 ZN A2 net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4 net_1 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6 net_2 B net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7 VDD C net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
M_i_1_1 net_0_0 A2 VSS VPW nfet_05v0 W=7.8e-07 L=6e-07
M_i_0_1 ZN A1 net_0_0 VPW nfet_05v0 W=7.8e-07 L=6e-07
M_i_0_0 net_0_1 A1 ZN VPW nfet_05v0 W=7.8e-07 L=6e-07
M_i_1_0 VSS A2 net_0_1 VPW nfet_05v0 W=7.8e-07 L=6e-07
M_i_2_0 ZN B VSS VPW nfet_05v0 W=5.15e-07 L=6e-07
M_i_3_0 VSS C ZN VPW nfet_05v0 W=5.15e-07 L=6e-07
M_i_3_1 ZN C VSS VPW nfet_05v0 W=5.15e-07 L=6e-07
M_i_2_1 VSS B ZN VPW nfet_05v0 W=5.15e-07 L=6e-07
M_i_5_1 ZN A2 net_1 VNW pfet_05v0 W=1.14e-06 L=5e-07
M_i_4_1 net_1 A1 ZN VNW pfet_05v0 W=1.14e-06 L=5e-07
M_i_4_0 ZN A1 net_1 VNW pfet_05v0 W=1.14e-06 L=5e-07
M_i_5_0 net_1 A2 ZN VNW pfet_05v0 W=1.14e-06 L=5e-07
M_i_6_0 net_2_0 B net_1 VNW pfet_05v0 W=1.14e-06 L=5e-07
M_i_7_0 VDD C net_2_0 VNW pfet_05v0 W=1.14e-06 L=5e-07
M_i_7_1 net_2_1 C VDD VNW pfet_05v0 W=1.14e-06 L=5e-07
M_i_6_1 net_1 B net_2_1 VNW pfet_05v0 W=1.14e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
M_i_1_3 net_0_0 A2 VSS VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_0_3 ZN A1 net_0_0 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_0_2 net_0_1 A1 ZN VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_1_2 VSS A2 net_0_1 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_1_1 net_0_2 A2 VSS VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_0_1 ZN A1 net_0_2 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_0_0 net_0_3 A1 ZN VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_1_0 VSS A2 net_0_3 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_2_0 ZN B VSS VPW nfet_05v0 W=4.6e-07 L=6e-07
M_i_3_0 VSS C ZN VPW nfet_05v0 W=4.6e-07 L=6e-07
M_i_3_1 ZN C VSS VPW nfet_05v0 W=4.6e-07 L=6e-07
M_i_2_1 VSS B ZN VPW nfet_05v0 W=4.6e-07 L=6e-07
M_i_2_2 ZN B VSS VPW nfet_05v0 W=4.6e-07 L=6e-07
M_i_3_2 VSS C ZN VPW nfet_05v0 W=4.6e-07 L=6e-07
M_i_3_3 ZN C VSS VPW nfet_05v0 W=4.6e-07 L=6e-07
M_i_2_3 VSS B ZN VPW nfet_05v0 W=4.6e-07 L=6e-07
M_i_5_3 ZN A2 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_3 net_1 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_2 ZN A1 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_2 net_1 A2 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_1 ZN A2 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_1 net_1 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_0 ZN A1 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_0 net_1 A2 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0 net_2_0 B net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 VDD C net_2_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 net_2_1 C VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_1 net_1 B net_2_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_2 net_2_2 B net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_2 VDD C net_2_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_3 net_2_3 C VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_3 net_1 B net_2_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
M_i_4 net_1 B2 VSS VPW nfet_05v0 W=7.1e-07 L=6e-07
M_i_3 ZN B1 net_1 VPW nfet_05v0 W=7.1e-07 L=6e-07
M_i_2 VSS C ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_1 net_0 A2 VSS VPW nfet_05v0 W=7.1e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=7.1e-07 L=6e-07
M_i_9 VDD B2 net_3 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_8 net_3 B1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7 net_2 C net_3 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6 ZN A2 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5 net_2 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
M_i_2_1 VSS C ZN VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_4_1 net_1_0 B2 VSS VPW nfet_05v0 W=7.15e-07 L=6e-07
M_i_3_1 ZN B1 net_1_0 VPW nfet_05v0 W=7.15e-07 L=6e-07
M_i_3_0 net_1_1 B1 ZN VPW nfet_05v0 W=7.15e-07 L=6e-07
M_i_4_0 VSS B2 net_1_1 VPW nfet_05v0 W=7.15e-07 L=6e-07
M_i_2_0 ZN C VSS VPW nfet_05v0 W=5.75e-07 L=6e-07
M_i_0_1 net_0_0 A1 ZN VPW nfet_05v0 W=7.15e-07 L=6e-07
M_i_1_1 VSS A2 net_0_0 VPW nfet_05v0 W=7.15e-07 L=6e-07
M_i_1_0 net_0_1 A2 VSS VPW nfet_05v0 W=7.15e-07 L=6e-07
M_i_0_0 ZN A1 net_0_1 VPW nfet_05v0 W=7.15e-07 L=6e-07
M_i_7_1 net_3 C net_2 VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_9_1 VDD B2 net_3 VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_8_1 net_3 B1 VDD VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_8_0 VDD B1 net_3 VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_9_0 net_3 B2 VDD VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_7_0 net_2 C net_3 VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_5_1 ZN A1 net_2 VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_6_1 net_2 A2 ZN VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_6_0 ZN A2 net_2 VNW pfet_05v0 W=1.12e-06 L=5e-07
M_i_5_0 net_2 A1 ZN VNW pfet_05v0 W=1.12e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
M_i_3_3 net_1_0 B1 ZN VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_4_3 VSS B2 net_1_0 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_4_2 net_1_1 B2 VSS VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_3_2 ZN B1 net_1_1 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_3_1 net_1_2 B1 ZN VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_4_1 VSS B2 net_1_2 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_4_0 net_1_3 B2 VSS VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_3_0 ZN B1 net_1_3 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_2_3 VSS C ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_2_2 ZN C VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_2_1 VSS C ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_2_0 ZN C VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_3 net_0_0 A1 ZN VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_1_3 VSS A2 net_0_0 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_1_2 net_0_1 A2 VSS VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_0_2 ZN A1 net_0_1 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_0_1 net_0_2 A1 ZN VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_1_1 VSS A2 net_0_2 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_1_0 net_0_3 A2 VSS VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_0_0 ZN A1 net_0_3 VPW nfet_05v0 W=7.7e-07 L=6e-07
M_i_8_3 net_3 B1 VDD VNW pfet_05v0 W=1.035e-06 L=5e-07
M_i_9_3 VDD B2 net_3 VNW pfet_05v0 W=1.035e-06 L=5e-07
M_i_9_2 net_3 B2 VDD VNW pfet_05v0 W=1.035e-06 L=5e-07
M_i_8_2 VDD B1 net_3 VNW pfet_05v0 W=1.035e-06 L=5e-07
M_i_8_1 net_3 B1 VDD VNW pfet_05v0 W=1.035e-06 L=5e-07
M_i_9_1 VDD B2 net_3 VNW pfet_05v0 W=1.035e-06 L=5e-07
M_i_9_0 net_3 B2 VDD VNW pfet_05v0 W=1.035e-06 L=5e-07
M_i_8_0 VDD B1 net_3 VNW pfet_05v0 W=1.035e-06 L=5e-07
M_i_7_3 net_3 C net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7_2 net_2 C net_3 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7_1 net_3 C net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7_0 net_2 C net_3 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_3 ZN A1 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_3 net_2 A2 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_2 ZN A2 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_2 net_2 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_1 ZN A1 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_1 net_2 A2 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_0 ZN A2 net_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_0 net_2 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
M_i_5 net_2 C2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4 ZN C1 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_1 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VSS B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 net_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_11 net_4 C2 VDD VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_10 VDD C1 net_4 VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_8 net_4 B1 net_3 VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_9 net_3 B2 net_4 VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_7 ZN A2 net_3 VNW pfet_05v0 W=1.16e-06 L=5e-07
M_i_6 net_3 A1 ZN VNW pfet_05v0 W=1.16e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
M_i_4_1 net_2_1 C1 ZN VPW nfet_05v0 W=8e-07 L=6e-07
M_i_5_1 VSS C2 net_2_1 VPW nfet_05v0 W=8e-07 L=6e-07
M_i_5_0 net_2_0 C2 VSS VPW nfet_05v0 W=8e-07 L=6e-07
M_i_4_0 ZN C1 net_2_0 VPW nfet_05v0 W=8e-07 L=6e-07
M_i_2_0 net_1_1 B1 ZN VPW nfet_05v0 W=8e-07 L=6e-07
M_i_3_0 VSS B2 net_1_1 VPW nfet_05v0 W=8e-07 L=6e-07
M_i_3_1 net_1_0 B2 VSS VPW nfet_05v0 W=8e-07 L=6e-07
M_i_2_1 ZN B1 net_1_0 VPW nfet_05v0 W=8e-07 L=6e-07
M_i_0_0 net_0_1 A1 ZN VPW nfet_05v0 W=8e-07 L=6e-07
M_i_1_0 VSS A2 net_0_1 VPW nfet_05v0 W=8e-07 L=6e-07
M_i_1_1 net_0_0 A2 VSS VPW nfet_05v0 W=8e-07 L=6e-07
M_i_0_1 ZN A1 net_0_0 VPW nfet_05v0 W=8e-07 L=6e-07
M_i_10_1 net_4 C1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11_1 VDD C2 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11_0 net_4 C2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_10_0 VDD C1 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8_0 net_4 B1 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9_0 net_3 B2 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9_1 net_4 B2 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8_1 net_3 B1 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0 ZN A1 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 net_3 A2 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 ZN A2 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_1 net_3 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
M_i_4_3 net_2_3 C1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_3 VSS C2 net_2_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_2 net_2_2 C2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_2 ZN C1 net_2_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_1 net_2_1 C1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 VSS C2 net_2_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_0 net_2_0 C2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 ZN C1 net_2_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_1_3 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS B2 net_1_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_1_2 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 ZN B1 net_1_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_1_1 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 VSS B2 net_1_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_3 net_1_0 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 ZN B1 net_1_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0_3 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 VSS A2 net_0_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0_2 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 net_0_1 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 VSS A2 net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 net_0_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 ZN A1 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10_3 net_4 C1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11_3 VDD C2 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11_2 net_4 C2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_10_2 VDD C1 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_10_1 net_4 C1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11_1 VDD C2 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11_0 net_4 C2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_10_0 VDD C1 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8_0 net_4 B1 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9_0 net_3 B2 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9_1 net_4 B2 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8_1 net_3 B1 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8_2 net_4 B1 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9_2 net_3 B2 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9_3 net_4 B2 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8_3 net_3 B1 net_4 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0 ZN A1 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 net_3 A2 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 ZN A2 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_1 net_3 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_2 ZN A1 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_2 net_3 A2 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_3 ZN A2 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_3 net_3 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
M_i_2 VSS I Z_neg VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VDD I Z_neg VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
M_i_2 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
M_i_2 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_4 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_5 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_6 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_7 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_2 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_3 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_4 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_5 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_4 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_5 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_6 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_7 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_8 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_9 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_10 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_11 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_2 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_3 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_4 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_5 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_4 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_5 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_6 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_7 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_4 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_5 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_6 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_7 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_8 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_9 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_10 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_11 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_12 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_13 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_14 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_15 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_2 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_3 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_4 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_5 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_6 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_7 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_12 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_13 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_14 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_15 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_4 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_5 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_6 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_7 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_8 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_9 VSS I Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_4 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_5 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_6 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_7 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_8 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_9 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_10 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_11 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_12 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_13 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_14 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_15 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_16 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_17 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_18 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_19 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_2 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_3 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_4 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_5 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_6 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_7 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_8 Z_neg I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_9 VDD I Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_12 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_13 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_14 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_15 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_16 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_17 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_18 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_19 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__bufz_1 EN I Z VDD VNW VPW VSS
M_XX27 VSS EN NEN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_XX44 VSS NEN NI_N VPW nfet_05v0 W=3.6e-07 L=6e-07
M_XX36 NI_N EN NI_P VPW nfet_05v0 W=3.6e-07 L=6e-07
M_XX43 NI_N I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_XX22 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX28 VDD EN NEN VNW pfet_05v0 W=6.2e-07 L=5e-07
M_XX45 NI_P EN VDD VNW pfet_05v0 W=6.2e-07 L=5e-07
M_XX39 NI_N NEN NI_P VNW pfet_05v0 W=6.2e-07 L=5e-07
M_XX46 NI_P I VDD VNW pfet_05v0 W=6.2e-07 L=5e-07
M_XX21 VDD NI_P Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__bufz_2 EN I Z VDD VNW VPW VSS
M_XX27 VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX44 VSS NEN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX36 NI_N EN NI_P VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX43 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22_4 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX28 VDD EN NEN VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX45 NI_P EN VDD VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX39 NI_N NEN NI_P VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX46 NI_P I VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX21 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX21_5 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__bufz_3 EN I Z VDD VNW VPW VSS
M_XX27 VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX44 VSS NEN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX36 NI_N EN NI_P VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX43 NI_N I VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_XX43_17 NI_N I VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_XX22 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22_4 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22_4_97 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX28 VDD EN NEN VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX45 NI_P EN VDD VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX39 NI_N NEN NI_P VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX46 NI_P I VDD VNW pfet_05v0 W=1.01e-06 L=5e-07
M_XX46_9 NI_P I VDD VNW pfet_05v0 W=1.01e-06 L=5e-07
M_XX21 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX21_5 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX21_5_72 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__bufz_4 EN I Z VDD VNW VPW VSS
M_XX27 VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX44 VSS NEN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX36 NI_N EN NI_P VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX43 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX43_17 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22_4 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22_4_97 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22_4_97_16 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX28 VDD EN NEN VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX45 NI_P EN VDD VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX39 NI_N NEN NI_P VNW pfet_05v0 W=9.45e-07 L=5e-07
M_XX46 NI_P I VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX46_9 NI_P I VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX21 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX21_5 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX21_5_72 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_XX21_5_72_5 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__bufz_8 EN I Z VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_34 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_88 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_33 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_99 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=9.45e-07 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=9.45e-07 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=9.45e-07 L=5e-07
M_mp14 NI_P I VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp14_10 VDD I NI_P VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp14_11 NI_P I VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp14_10_8 VDD I NI_P VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57_75 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56_111 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_106 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_58 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__bufz_12 EN I Z VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10_0 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17_30 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_34 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_88 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_33 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_99 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_35 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_80 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_34 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_89 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=9.45e-07 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=9.45e-07 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=9.45e-07 L=5e-07
M_mp14 NI_P I VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp14_10 VDD I NI_P VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp14_11 NI_P I VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp14_10_8 VDD I NI_P VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp14_11_21 NI_P I VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp14_10_8_17 VDD I NI_P VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57_75 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56_111 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_106 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_58 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57_69 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56_105 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_96 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_57 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__bufz_16 EN I Z VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn17 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_34 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_41 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10_30 NI_N I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17_61 VSS I NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_34 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_88 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_33 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_99 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_34_75 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_88_82 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_33_198 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_99_125 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_137 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_181 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_65 Z NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_118 VSS NI_N Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=9.2e-07 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=9.2e-07 L=5e-07
M_mp14 NI_P I VDD VNW pfet_05v0 W=1.15e-06 L=5e-07
M_mp14_10 VDD I NI_P VNW pfet_05v0 W=1.15e-06 L=5e-07
M_mp14_11 NI_P I VDD VNW pfet_05v0 W=1.15e-06 L=5e-07
M_mp14_10_8 VDD I NI_P VNW pfet_05v0 W=1.15e-06 L=5e-07
M_mp14_7 NI_P I VDD VNW pfet_05v0 W=1.15e-06 L=5e-07
M_mp14_10_32 VDD I NI_P VNW pfet_05v0 W=1.15e-06 L=5e-07
M_mp14_11_55 NI_P I VDD VNW pfet_05v0 W=1.15e-06 L=5e-07
M_mp14_10_8_20 VDD I NI_P VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57_75 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56_111 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_106 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_58 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57_75_85 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56_111_134 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_106_111 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_58_95 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_57_97 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_56_133 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_12_126 Z NI_P VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
M_mp4_153 VDD NI_P Z VNW pfet_05v0 W=1.175e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
M_i_2 VSS I Z_neg VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=4.95e-07 L=6e-07
M_i_3 VDD I Z_neg VNW pfet_05v0 W=5.25e-07 L=5e-07
M_i_3_0 VDD I Z_neg VNW pfet_05v0 W=5.25e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
M_i_2 VSS I Z_neg VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_3 VDD I Z_neg VNW pfet_05v0 W=1.02e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=6.05e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=4.55e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=4.55e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=4.55e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=4.55e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=12.2e-07 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=12.2e-07 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=12.2e-07 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=12.2e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=6.05e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=4.55e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=4.55e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=4.55e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=4.55e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_2_2 Z_neg I VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=4.3e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=4.3e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=4.3e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=4.3e-07 L=6e-07
M_i_0_4 Z Z_neg VSS VPW nfet_05v0 W=4.3e-07 L=6e-07
M_i_0_5 VSS Z_neg Z VPW nfet_05v0 W=4.3e-07 L=6e-07
M_i_0_6 Z Z_neg VSS VPW nfet_05v0 W=4.3e-07 L=6e-07
M_i_0_7 VSS Z_neg Z VPW nfet_05v0 W=4.3e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_2 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_3 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_2 Z_neg I VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_3 VSS I Z_neg VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_4 Z_neg I VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_4 Z Z_neg VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_5 VSS Z_neg Z VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_6 Z Z_neg VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_7 VSS Z_neg Z VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_8 Z Z_neg VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_9 VSS Z_neg Z VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_10 Z Z_neg VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_11 VSS Z_neg Z VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_2 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_3 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_4 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_5 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_2_2 Z_neg I VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_2_3 VSS I Z_neg VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_2_4 Z_neg I VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_2_5 VSS I Z_neg VPW nfet_05v0 W=4.05e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_4 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_5 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_6 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_7 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_8 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_9 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_10 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_11 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_12 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_13 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_14 Z Z_neg VSS VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_0_15 VSS Z_neg Z VPW nfet_05v0 W=4.85e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_2 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_3 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_4 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_5 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_6 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_7 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_12 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_13 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_14 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_15 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_2_1 VSS I Z_neg VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_2_2 Z_neg I VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_2_3 VSS I Z_neg VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_2_4 Z_neg I VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_2_5 VSS I Z_neg VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_2_6 Z_neg I VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_2_7 VSS I Z_neg VPW nfet_05v0 W=3.8e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_4 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_5 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_6 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_7 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_8 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_9 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_10 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_11 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_12 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_13 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_14 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_15 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_16 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_17 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_18 Z Z_neg VSS VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_0_19 VSS Z_neg Z VPW nfet_05v0 W=4.7e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_1 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_2 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_3 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_4 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_5 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_6 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_7 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_8 Z_neg I VDD VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_3_9 VDD I Z_neg VNW pfet_05v0 W=0.82e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_12 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_13 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_14 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_15 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_16 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_17 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_18 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_19 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
M_i_0 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_1 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_3 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VNW VPW VSS
M_i_0_0_x8_0 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_0_x8_1 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_0_x8_2 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_0_x8_3 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_0_x8_4 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_0_x8_5 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_0_x8_6 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_0_x8_7 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_1_0_x8_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_4 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_5 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_6 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_7 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_3 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_4 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_5 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_6 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_7 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_8 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_9 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_10 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_11 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkinv_16 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_3 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_4 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_5 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_6 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_7 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_8 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_9 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_10 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_11 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_12 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_13 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_14 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_15 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_12 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_13 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_14 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_15 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__clkinv_20 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_3 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_4 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_5 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_6 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_7 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_8 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_9 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_10 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_11 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_12 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_13 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_14 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_15 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_16 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_17 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_18 ZN I VSS VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_0_19 VSS I ZN VPW nfet_05v0 W=4.8e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_12 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_13 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_14 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_15 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_16 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_17 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_18 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_19 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VNW VPW VSS
M_tn9 ncki CLKN VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn16 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 VSS D net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net2 cki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net5 ncki net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 VSS net10 net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 net5 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 ncki net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net7 cki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 VSS net1 net7 VPW nfet_05v0 W=6.3e-07 L=6e-07
M_tn5 net1 net0 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_tn6 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp9 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp16 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp10 VDD D net2 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp11 net5 ncki net2 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp0 net4 cki net5 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp1 VDD net10 net4 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp15 net10 net5 VDD VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp7 net0 cki net10 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp6 net7 ncki net0 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp2 VDD net1 net7 VNW pfet_05v0 W=1.075e-06 L=5e-07
M_tp3 net1 net0 VDD VNW pfet_05v0 W=1.075e-06 L=5e-07
M_tp4 Q net1 VDD VNW pfet_05v0 W=11.3e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnq_2 D CLKN Q VDD VNW VPW VSS
M_tn9 ncki CLKN VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn16 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 VSS D net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net2 cki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net5 ncki net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 VSS net10 net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 net5 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 ncki net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net7 cki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 VSS net1 net7 VPW nfet_05v0 W=9.45e-07 L=6e-07
M_tn5 net1 net0 VSS VPW nfet_05v0 W=9.45e-07 L=6e-07
M_tn6_7 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp9 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp16 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp10 VDD D net2 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp11 net5 ncki net2 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp0 net4 cki net5 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp1 VDD net10 net4 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp15 net10 net5 VDD VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp7 net0 cki net10 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp6 net7 ncki net0 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp2 VDD net1 net7 VNW pfet_05v0 W=1.075e-06 L=5e-07
M_tp3 net1 net0 VDD VNW pfet_05v0 W=1.075e-06 L=5e-07
M_tp4_13 Q net1 VDD VNW pfet_05v0 W=10.95e-07 L=5e-07
M_tp4 Q net1 VDD VNW pfet_05v0 W=10.95e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnq_4 D CLKN Q VDD VNW VPW VSS
M_tn9 ncki CLKN VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn16 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 VSS D net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net2 cki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net5 ncki net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 VSS net10 net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 net5 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 ncki net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net7 cki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 VSS net1 net7 VPW nfet_05v0 W=9.45e-07 L=6e-07
M_tn5 net1 net0 VSS VPW nfet_05v0 W=9.45e-07 L=6e-07
M_tn6_7 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6_7_61 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6_49 Q net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp9 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp16 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp10 VDD D net2 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp11 net5 ncki net2 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp0 net4 cki net5 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp1 VDD net10 net4 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp15 net10 net5 VDD VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp7 net0 cki net10 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp6 net7 ncki net0 VNW pfet_05v0 W=4.95e-07 L=5e-07
M_tp2 VDD net1 net7 VNW pfet_05v0 W=1.075e-06 L=5e-07
M_tp3 net1 net0 VDD VNW pfet_05v0 W=1.075e-06 L=5e-07
M_tp4_13 Q net1 VDD VNW pfet_05v0 W=10.95e-07 L=5e-07
M_tp4 Q net1 VDD VNW pfet_05v0 W=10.95e-07 L=5e-07
M_tp4_13_64 Q net1 VDD VNW pfet_05v0 W=10.95e-07 L=5e-07
M_tp4_55 Q net1 VDD VNW pfet_05v0 W=10.95e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VNW VPW VSS
M_tn13 ncki CLKN VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn10 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn11 net6 D VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn15 net6 cki net1 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn14 net1 ncki net15 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn0 net8 ncki net2 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn1 net11 cki net8 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=4e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=7.95e-07 L=6e-07
M_tp11 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp8 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp9 VDD D net6 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp15 net1 ncki net6 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp7 net9 cki net1 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp2 net2 cki net8 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net8 ncki net11 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=0.94e-06 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=0.94e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.175e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2 D RN CLKN Q VDD VNW VPW VSS
M_tn13 ncki CLKN VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn10 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn11 net6 D VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn15 net6 cki net1 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn14 net1 ncki net15 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn0 net8 ncki net2 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn1 net11 cki net8 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=8.25e-07 L=6e-07
M_tn3_42 Q net4 VSS VPW nfet_05v0 W=7.95e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=7.95e-07 L=6e-07
M_tp11 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp8 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp9 VDD D net6 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp15 net1 ncki net6 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp7 net9 cki net1 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp2 net2 cki net8 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net8 ncki net11 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=1.09e-06 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=1.09e-06 L=5e-07
M_tp1_40 Q net4 VDD VNW pfet_05v0 W=1.185e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.185e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4 D RN CLKN Q VDD VNW VPW VSS
M_tn13 ncki CLKN VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn10 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn11 net6 D VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn15 net6 cki net1 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn14 net1 ncki net15 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn0 net8 ncki net2 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn1 net11 cki net8 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=8.25e-07 L=6e-07
M_tn3_42 Q net4 VSS VPW nfet_05v0 W=7.95e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=7.95e-07 L=6e-07
M_tn3_42_63 Q net4 VSS VPW nfet_05v0 W=7.95e-07 L=6e-07
M_tn3_69 Q net4 VSS VPW nfet_05v0 W=7.95e-07 L=6e-07
M_tp11 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp8 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp9 VDD D net6 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp15 net1 ncki net6 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp7 net9 cki net1 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=7.6e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp2 net2 cki net8 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net8 ncki net11 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_tp1_40 Q net4 VDD VNW pfet_05v0 W=1.205e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.205e-06 L=5e-07
M_tp1_40_64 Q net4 VDD VNW pfet_05v0 W=1.205e-06 L=5e-07
M_tp1_66 Q net4 VDD VNW pfet_05v0 W=1.205e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1 D RN SETN CLKN Q VDD VNW VPW VSS
M_tn2 ncki CLKN VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn1 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 net14 D VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn8 net14 cki net3 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn5 net3 ncki net16 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net5 ncki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net7 cki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp2 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp1 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 VDD D net14 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp10 net3 ncki net14 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp7 net13 cki net3 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=8.05e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=8.05e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp20 net4 cki net5 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp19 net5 ncki net7 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2 D RN SETN CLKN Q VDD VNW VPW VSS
M_tn2 ncki CLKN VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn1 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 net14 D VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn8 net14 cki net3 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn5 net3 ncki net16 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net5 ncki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net7 cki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn19_16 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp2 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp1 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 VDD D net14 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp10 net3 ncki net14 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp7 net13 cki net3 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=8.05e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=8.05e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp20 net4 cki net5 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp19 net5 ncki net7 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp17_9 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4 D RN SETN CLKN Q VDD VNW VPW VSS
M_tn2 ncki CLKN VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn1 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 net14 D VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn8 net14 cki net3 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn5 net3 ncki net16 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net5 ncki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net7 cki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn19_16 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn19_16_44 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn19_64 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp2 ncki CLKN VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp1 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 VDD D net14 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp10 net3 ncki net14 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp7 net13 cki net3 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=4.1e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=8.05e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=8.05e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp20 net4 cki net5 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp19 net5 ncki net7 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=8.75e-07 L=5e-07
M_tp17_9 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp17_9_60 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp17_57 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VNW VPW VSS
M_tn0 ncki CLKN VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn3 cki ncki VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn10 net13 D VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn6 net13 cki net3 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn4 net3 ncki net14 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn13 net5 ncki net4 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn12 net7 cki net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=4.35e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=3.1e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=3.75e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp0 ncki CLKN VDD VNW pfet_05v0 W=9.4e-07 L=5e-07
M_tp4 cki ncki VDD VNW pfet_05v0 W=9.4e-07 L=5e-07
M_tp8 VDD D net13 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp9 net3 ncki net13 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp6 net10 cki net3 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=5.7e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp18 net5 cki net4 VNW pfet_05v0 W=5.35e-07 L=5e-07
M_tp17 net7 ncki net5 VNW pfet_05v0 W=6.5e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=7.05e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=5.8e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=6.55e-07 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2 D SETN CLKN Q VDD VNW VPW VSS
M_tn0 ncki CLKN VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn3 cki ncki VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn10 net13 D VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn6 net13 cki net3 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn4 net3 ncki net14 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn13 net5 ncki net4 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn12 net7 cki net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=4.35e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=3.1e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=3.75e-07 L=6e-07
M_tn16_30 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp0 ncki CLKN VDD VNW pfet_05v0 W=9.4e-07 L=5e-07
M_tp4 cki ncki VDD VNW pfet_05v0 W=9.4e-07 L=5e-07
M_tp8 VDD D net13 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp9 net3 ncki net13 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp6 net10 cki net3 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=5.7e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp18 net5 cki net4 VNW pfet_05v0 W=5.35e-07 L=5e-07
M_tp17 net7 ncki net5 VNW pfet_05v0 W=6.5e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=7.05e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=5.8e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=6.55e-07 L=5e-07
M_tp14_24 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4 D SETN CLKN Q VDD VNW VPW VSS
M_tn0 ncki CLKN VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn3 cki ncki VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn10 net13 D VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn6 net13 cki net3 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn4 net3 ncki net14 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn13 net5 ncki net4 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn12 net7 cki net5 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=4.35e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=3.1e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=3.75e-07 L=6e-07
M_tn16_30 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_30_46 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_51 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp0 ncki CLKN VDD VNW pfet_05v0 W=9.4e-07 L=5e-07
M_tp4 cki ncki VDD VNW pfet_05v0 W=9.4e-07 L=5e-07
M_tp8 VDD D net13 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp9 net3 ncki net13 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp6 net10 cki net3 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=6.05e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=5.7e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp18 net5 cki net4 VNW pfet_05v0 W=5.35e-07 L=5e-07
M_tp17 net7 ncki net5 VNW pfet_05v0 W=6.5e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=7.05e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=5.8e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=6.55e-07 L=5e-07
M_tp14_24 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp14_24_63 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp14_44 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
M_tn3 VSS CLK ncki VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn4 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn5 net5 ncki VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net4 D net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net6 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS net0 net6 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net0 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 net2 cki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net1 ncki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 VSS net3 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 net3 net2 VSS VPW nfet_05v0 W=4e-07 L=6e-07
M_tn1 Q net3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp3 VDD CLK ncki VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp4 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp12 net7 cki VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp11 net4 D net7 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp6 net8 ncki net4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp5 VDD net0 net8 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp0 net0 net4 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp7 net2 ncki net0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp9 net1x cki net2 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp10 VDD net3 net1x VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp8 net3 net2 VDD VNW pfet_05v0 W=8e-07 L=5e-07
M_tp1 Q net3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
M_tn3 VSS CLK ncki VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn4 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn5 net5 ncki VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net4 D net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net6 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS net0 net6 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net0 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 net2 cki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net1 ncki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 VSS net3 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 net3 net2 VSS VPW nfet_05v0 W=4e-07 L=6e-07
M_tn1 Q net3 VSS VPW nfet_05v0 W=1.64e-06 L=6e-07
M_tp3 VDD CLK ncki VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp4 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp12 net7 cki VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp11 net4 D net7 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp6 net8 ncki net4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp5 VDD net0 net8 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp0 net0 net4 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp7 net2 ncki net0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp9 net1x cki net2 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp10 VDD net3 net1x VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp8 net3 net2 VDD VNW pfet_05v0 W=8e-07 L=5e-07
M_tp1 Q net3 VDD VNW pfet_05v0 W=2.44e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
M_tn3 VSS CLK ncki VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn4 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn5 net5 ncki VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net4 D net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net6 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS net0 net6 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net0 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 net2 cki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net1 ncki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 VSS net3 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 net3 net2 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn10_6 net3 net2 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn1_39 Q net3 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn1_18_47 Q net3 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn1 Q net3 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn1_18 Q net3 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp3 VDD CLK ncki VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp4 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp12 net7 cki VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp11 net4 D net7 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp6 net8 ncki net4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp5 VDD net0 net8 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp0 net0 net4 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp7 net2 ncki net0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp9 net1x cki net2 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp10 VDD net3 net1x VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp8 net3 net2 VDD VNW pfet_05v0 W=9.45e-07 L=5e-07
M_tp8_10 net3 net2 VDD VNW pfet_05v0 W=9.45e-07 L=5e-07
M_tp1_58 Q net3 VDD VNW pfet_05v0 W=12.2e-07 L=5e-07
M_tp1_16_34 Q net3 VDD VNW pfet_05v0 W=12.2e-07 L=5e-07
M_tp1 Q net3 VDD VNW pfet_05v0 W=12.2e-07 L=5e-07
M_tp1_16 Q net3 VDD VNW pfet_05v0 W=12.2e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
M_tn10 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn13 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn11 net10 D VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 ncki net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 cki net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net8 cki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net11 ncki net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=4e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp8 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp11 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp9 VDD D net10 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp15 net1 cki net10 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp7 net9 ncki net1 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp2 net2 ncki net8 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net8 cki net11 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=1e-06 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=1e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VNW VPW VSS
M_tn10 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn13 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn11 net10 D VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 ncki net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 cki net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net8 cki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net11 ncki net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn3_15 Q net4 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp8 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp11 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp9 VDD D net10 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp15 net1 cki net10 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp7 net9 ncki net1 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp2 net2 ncki net8 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net8 cki net11 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1_13 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VNW VPW VSS
M_tn10 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn13 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn11 net10 D VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 ncki net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 cki net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net8 cki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net11 ncki net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn3_15 Q net4 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn3_15_13 Q net4 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn3_10 Q net4 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp8 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp11 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp9 VDD D net10 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp15 net1 cki net10 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp7 net9 ncki net1 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp2 net2 ncki net8 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net8 cki net11 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1_13 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1_13_25 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1_30 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 D RN SETN CLK Q VDD VNW VPW VSS
M_tn1 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn2 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 net14 D VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn8 net14 ncki net3 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn5 net3 cki net16 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn14 net5 cki net4 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn13 net7 ncki net5 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp1 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp2 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 VDD D net14 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp10 net3 cki net14 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp7 net13 ncki net3 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=7.55e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=7.55e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp20 net4 ncki net5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp19 net5 cki net7 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2 D RN SETN CLK Q VDD VNW VPW VSS
M_tn1 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn2 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 net14 D VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn8 net14 ncki net3 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn5 net3 cki net16 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn14 net5 cki net4 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn13 net7 ncki net5 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn19_39 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp1 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp2 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 VDD D net14 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp10 net3 cki net14 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp7 net13 ncki net3 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=3.65e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=7.55e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=7.55e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp20 net4 ncki net5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp19 net5 cki net7 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp17_33 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4 D RN SETN CLK Q VDD VNW VPW VSS
M_tn1 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn2 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 net14 D VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn8 net14 ncki net3 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn5 net3 cki net16 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn14 net5 cki net4 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn13 net7 ncki net5 VPW nfet_05v0 W=5.05e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn19_39 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn19_39_20 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn19_24 Q net6 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp1 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp2 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 VDD D net14 VNW pfet_05v0 W=4.75e-07 L=5e-07
M_tp10 net3 cki net14 VNW pfet_05v0 W=4.75e-07 L=5e-07
M_tp7 net13 ncki net3 VNW pfet_05v0 W=4.75e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=4.75e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=6.9e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=6.9e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp20 net4 ncki net5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp19 net5 cki net7 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=7.7e-07 L=5e-07
M_tp17_33 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp17_33_0 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp17_16 Q net6 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VNW VPW VSS
M_tn3 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn10 net13 D VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net13 ncki net3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net3 cki net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp4 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp8 VDD D net13 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp9 net3 cki net13 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp6 net10 ncki net3 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=5.85e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=5.85e-07 L=5e-07
M_tp18 net5 ncki net4 VNW pfet_05v0 W=4.15e-07 L=5e-07
M_tp17 net7 cki net5 VNW pfet_05v0 W=4.15e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VNW VPW VSS
M_tn3 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn10 net13 D VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net13 ncki net3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net3 cki net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_7 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp4 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp8 VDD D net13 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp9 net3 cki net13 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp6 net10 ncki net3 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=5.85e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=5.85e-07 L=5e-07
M_tp18 net5 ncki net4 VNW pfet_05v0 W=4.15e-07 L=5e-07
M_tp17 net7 cki net5 VNW pfet_05v0 W=4.15e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=1.055e-06 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp14_2 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VNW VPW VSS
M_tn3 ncki CLK VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn0 cki ncki VSS VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn10 net13 D VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net13 ncki net3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net3 cki net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=4.05e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn18_45 net6 net5 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_7 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_23 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_7_36 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp4 ncki CLK VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp0 cki ncki VDD VNW pfet_05v0 W=8.65e-07 L=5e-07
M_tp8 VDD D net13 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp9 net3 cki net13 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp6 net10 ncki net3 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=5.05e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=5.85e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=5.85e-07 L=5e-07
M_tp18 net5 ncki net4 VNW pfet_05v0 W=4.15e-07 L=5e-07
M_tp17 net7 cki net5 VNW pfet_05v0 W=4.15e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=1.055e-06 L=5e-07
M_tp16_52 net6 net5 VDD VNW pfet_05v0 W=1.055e-06 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp14_2 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp14_19 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp14_2_27 VDD net6 Q VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlya_1 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 VSS Z_neg net_2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_6 net_3 net_2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 VDD Z_neg net_2 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_3 net_2 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 VSS Z_neg net_2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_6 net_3 net_2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 VDD Z_neg net_2 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_3 net_2 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlya_4 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 VSS Z_neg net_2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_6 net_3 net_2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_2 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1_15 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 VDD Z_neg net_2 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_3 net_2 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_34 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14_19 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_2 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_2 net_6 VPW nfet_05v0 W=3.65e-07 L=0.600000U
M_i_3_6 net_6 net_2 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_2 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_2 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_2 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyb_2 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_2 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_2 net_6 VPW nfet_05v0 W=3.65e-07 L=0.600000U
M_i_3_6 net_6 net_2 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_2 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_2 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_2 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyb_4 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_2 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_2 net_6 VPW nfet_05v0 W=3.65e-07 L=0.600000U
M_i_3_6 net_6 net_2 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_2 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1_15 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_2 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_2 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_2 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_34 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14_19 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_7 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26 net_9 net_7 net_13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30 net_13 net_7 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_1 net_8 net_9 net_11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4 net_11 net_9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_8 net_6 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3_6 net_6 net_8 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_7 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35 net_12 net_7 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47 net_9 net_7 net_12 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9 net_10 net_9 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22 net_8 net_9 net_10 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_8 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_8 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyc_2 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_7 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26 net_9 net_7 net_13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30 net_13 net_7 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_1 net_8 net_9 net_11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4 net_11 net_9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_8 net_6 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3_6 net_6 net_8 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_2 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_7 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35 net_12 net_7 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47 net_9 net_7 net_12 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9 net_10 net_9 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22 net_8 net_9 net_10 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_8 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_8 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_16 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyc_4 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_7 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26 net_9 net_7 net_13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30 net_13 net_7 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_1 net_8 net_9 net_11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4 net_11 net_9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_8 net_6 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3_6 net_6 net_8 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_2 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_2_36 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_7 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35 net_12 net_7 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47 net_9 net_7 net_12 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9 net_10 net_9 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22 net_8 net_9 net_10 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_8 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_8 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_16 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_32 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_16_16 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_7 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26 net_9 net_7 net_13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30 net_13 net_7 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_1 net_15 net_9 net_11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4 net_11 net_9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26_13 net_16 net_15 net_18 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30_34 net_18 net_15 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_10 net_14 net_16 net_19 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4_49 net_19 net_16 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_14 net_6 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3_6 net_6 net_14 VSS VPW nfet_05v0  W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_7 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35 net_12 net_7 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47 net_9 net_7 net_12 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9 net_10 net_9 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22 net_15 net_9 net_10 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35_50 net_17 net_15 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47_46 net_16 net_15 net_17 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9_2 net_20 net_16 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22_38 net_14 net_16 net_20 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_14 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_14 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyd_2 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_7 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26 net_9 net_7 net_13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30 net_13 net_7 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_1 net_15 net_9 net_11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4 net_11 net_9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26_13 net_16 net_15 net_18 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30_34 net_18 net_15 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_10 net_14 net_16 net_19 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4_49 net_19 net_16 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_14 net_6 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3_6 net_6 net_14 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_7 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35 net_12 net_7 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47 net_9 net_7 net_12 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9 net_10 net_9 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22 net_15 net_9 net_10 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35_50 net_17 net_15 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47_46 net_16 net_15 net_17 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9_2 net_20 net_16 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22_38 net_14 net_16 net_20 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_14 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_14 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VNW VPW VSS
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_7 Z_neg net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 net_1 Z_neg VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26 net_9 net_7 net_13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30 net_13 net_7 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_1 net_15 net_9 net_11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4 net_11 net_9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_26_13 net_16 net_15 net_18 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_30_34 net_18 net_15 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0_10 net_14 net_16 net_19 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_4_49 net_19 net_16 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_21 net_3 net_14 net_6 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_3_6 net_6 net_14 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_2 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0_18_1_15 Z net_3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0 net_0 Z_neg VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1 net_7 Z_neg net_0 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35 net_12 net_7 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47 net_9 net_7 net_12 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9 net_10 net_9 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22 net_15 net_9 net_10 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_35_50 net_17 net_15 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_47_46 net_16 net_15 net_17 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_9_2 net_20 net_16 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_22_38 net_14 net_16 net_20 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_0_29 net_5 net_14 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_1_39 net_3 net_14 net_5 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_34 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0_0_14_19 Z net_3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__endcap VDD VNW VPW VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fill_4 VDD VNW VPW VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fill_8 VDD VNW VPW VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fill_16 VDD VNW VPW VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fill_32 VDD VNW VPW VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fill_64 VDD VNW VPW VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
M_i_17 net_1 net_0 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_19 VDD net_1 net_0 VNW pfet_05v0 W=1.22e-06 L=1e-06
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
M_i_17 net_3 net_2 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23 net_4 net_5 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_19 VDD net_3 net_2 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7 VDD net_4 net_5 VNW pfet_05v0 W=1.22e-06 L=1e-06
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
M_i_17 net_3 net_2 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23 net_4 net_5 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24 net_7 net_9 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55 net_6 net_8 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_19 VDD net_3 net_2 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7 VDD net_4 net_5 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33 VDD net_7 net_9 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23 VDD net_6 net_8 VNW pfet_05v0 W=1.22e-06 L=1e-06
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
M_i_17 net_3 net_2 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23 net_4 net_5 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24 net_7 net_9 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55 net_6 net_8 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_27 net_17 net_14 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_63 net_16 net_15 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24_22 net_13 net_11 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55_93 net_12 net_10 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_19 VDD net_3 net_2 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7 VDD net_4 net_5 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33 VDD net_7 net_9 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23 VDD net_6 net_8 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_94 VDD net_17 net_14 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_87 VDD net_16 net_15 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33_95 VDD net_13 net_11 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23_23 VDD net_12 net_10 VNW pfet_05v0 W=1.22e-06 L=1e-06
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
M_i_17 net_3 net_2 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23 net_4 net_5 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24 net_7 net_9 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55 net_6 net_8 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_27 net_17 net_14 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_63 net_16 net_15 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24_22 net_13 net_11 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55_93 net_12 net_10 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_20 net_30 net_26 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_59 net_25 net_20 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24_135 net_23 net_28 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55_90 net_33 net_18 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_27_139 net_31 net_29 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_63_82 net_32 net_24 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_24_22_30 net_22 net_27 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_17_23_55_93_110 net_19 net_21 VSS VPW nfet_05v0 W=8.2e-07 L=1e-06
M_i_19 VDD net_3 net_2 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7 VDD net_4 net_5 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33 VDD net_7 net_9 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23 VDD net_6 net_8 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_94 VDD net_17 net_14 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_87 VDD net_16 net_15 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33_95 VDD net_13 net_11 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23_23 VDD net_12 net_10 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_95 VDD net_30 net_26 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_188 VDD net_25 net_20 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33_98 VDD net_23 net_28 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23_16 VDD net_33 net_18 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_94_91 VDD net_31 net_29 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_87_65 VDD net_32 net_24 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_33_95_109 VDD net_22 net_27 VNW pfet_05v0 W=1.22e-06 L=1e-06
M_i_19_7_23_23_99 VDD net_19 net_21 VNW pfet_05v0 W=1.22e-06 L=1e-06
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__hold Z VDD VNW VPW VSS
M_MU11 Z net8 VSS VPW nfet_05v0 W=3.2e-07 L=2e-06
M_u3 VSS Z net8 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MU12 Z net8 VDD VNW pfet_05v0 W=3.2e-07 L=2e-06
M_u7 VDD Z net8 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__icgtn_1 CLKN E TE Q VDD VNW VPW VSS
M_MU19 VSS TE net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU20 net50 E VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU75_M_u2 Q d3 VSS VPW nfet_05v0 W=6.25e-07 L=6e-07
M_MI81 net58 TE VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU17 net61 E net58 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU81_M_u3 VDD CLKN CP VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MI1_M_u2 d3 CLKN XI1-net8 VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MU75_M_u3 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU82_M_u2 NCP CP VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU81_M_u2 VSS CLKN CP VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI1_M_u4 VSS CLKN d3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU16 net53 CP net61 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI90 net067 NCP net53 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI88 VDD QD net067 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MU82_M_u3 NCP CP VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI95_M_u3 VDD net53 QD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI1_M_u1 XI1-net8 net36 VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MI82 net53 NCP net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI91 net038 CP net53 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI92 VSS QD net038 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI95_M_u2 VSS net53 QD VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI89_M_u2 net36 QD VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI1_M_u3 d3 net36 VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI89_M_u3 net36 QD VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__icgtn_2 CLKN E TE Q VDD VNW VPW VSS
M_MU19 VSS TE net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU20 net50 E VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU75_M_u2 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU75_M_u2_19 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MI81 net58 TE VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU17 net61 E net58 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU81_M_u3 VDD CLKN CP VNW pfet_05v0 W=1.155e-06 L=5e-07
M_MI1_M_u2 d3 CLKN XI1-net8 VNW pfet_05v0 W=1.155e-06 L=5e-07
M_MU75_M_u3 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3_1 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU82_M_u2 NCP CP VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU81_M_u2 VSS CLKN CP VPW nfet_05v0 W=4.75e-07 L=6e-07
M_MI1_M_u4 VSS CLKN d3 VPW nfet_05v0 W=4.75e-07 L=6e-07
M_MU16 net53 CP net61 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI90 net067 NCP net53 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI88 VDD QD net067 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MU82_M_u3 NCP CP VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI95_M_u3 VDD net53 QD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI1_M_u1 XI1-net8 net36 VDD VNW pfet_05v0 W=1.155e-06 L=5e-07
M_MI82 net53 NCP net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI91 net038 CP net53 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI92 VSS QD net038 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI95_M_u2 VSS net53 QD VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI89_M_u2 net36 QD VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI1_M_u3 d3 net36 VSS VPW nfet_05v0 W=4.75e-07 L=6e-07
M_MI89_M_u3 net36 QD VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__icgtn_4 CLKN E TE Q VDD VNW VPW VSS
M_MU19 VSS TE net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU20 net50 E VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU75_M_u2 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU75_M_u2_19 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU75_M_u2_33 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU75_M_u2_19_5 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MI81 net58 TE VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU17 net61 E net58 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU81_M_u3 VDD CLKN CP VNW pfet_05v0 W=1.155e-06 L=5e-07
M_MI1_M_u2 d3 CLKN XI1-net8 VNW pfet_05v0 W=1.155e-06 L=5e-07
M_MU75_M_u3 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3_1 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3_2 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3_1_35 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU82_M_u2 NCP CP VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU81_M_u2 VSS CLKN CP VPW nfet_05v0 W=4.75e-07 L=6e-07
M_MI1_M_u4 VSS CLKN d3 VPW nfet_05v0 W=4.75e-07 L=6e-07
M_MU16 net53 CP net61 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI90 net067 NCP net53 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI88 VDD QD net067 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MU82_M_u3 NCP CP VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI95_M_u3 VDD net53 QD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI1_M_u1 XI1-net8 net36 VDD VNW pfet_05v0 W=1.155e-06 L=5e-07
M_MI82 net53 NCP net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI91 net038 CP net53 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI92 VSS QD net038 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI95_M_u2 VSS net53 QD VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI89_M_u2 net36 QD VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI1_M_u3 d3 net36 VSS VPW nfet_05v0 W=4.75e-07 L=6e-07
M_MI89_M_u3 net36 QD VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__icgtp_1 CLK E TE Q VDD VNW VPW VSS
M_MU19 net50 TE VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU20 VSS E net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU81_M_u2 NCK CLK VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_MU75_M_u2 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MI81 VDD TE net58 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU17 net58 E net61 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU82_M_u3 CK NCK VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MU81_M_u3 VDD CLK NCK VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MI85_M_u1 d3 CLK VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MU75_M_u3 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MI82 net50 NCK net53 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI91 net53 CK net033 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI92 net033 QD VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI80_M_u2 VSS net53 QD VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU82_M_u2 VSS NCK CK VPW nfet_05v0 W=3.9e-07 L=6e-07
M_MI85_M_u3 XI85-net6 CLK d3 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_MI85_M_u4 VSS QD XI85-net6 VPW nfet_05v0 W=3.9e-07 L=6e-07
M_MU16 net61 CK net53 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI90 net53 NCK net062 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI88 net062 QD VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI80_M_u3 VDD net53 QD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI85_M_u2 VDD QD d3 VNW pfet_05v0 W=9.2e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__icgtp_2 CLK E TE Q VDD VNW VPW VSS
M_MU19 net50 TE VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU20 VSS E net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU81_M_u2 NCK CLK VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_MU75_M_u2 Q d3 VSS VPW nfet_05v0 W=6.25e-07 L=6e-07
M_MU75_M_u2_22 Q d3 VSS VPW nfet_05v0 W=6.25e-07 L=6e-07
M_MI81 VDD TE net58 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU17 net58 E net61 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU82_M_u3 CK NCK VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MU81_M_u3 VDD CLK NCK VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MI85_M_u1 d3 CLK VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3_3 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MI82 net50 NCK net53 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI91 net53 CK net033 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI92 net033 QD VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI80_M_u2 VSS net53 QD VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU82_M_u2 VSS NCK CK VPW nfet_05v0 W=3.9e-07 L=6e-07
M_MI85_M_u3 XI85-net6 CLK d3 VPW nfet_05v0 W=6.25e-07 L=6e-07
M_MI85_M_u4 VSS QD XI85-net6 VPW nfet_05v0 W=6.25e-07 L=6e-07
M_MU16 net61 CK net53 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI90 net53 NCK net062 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI88 net062 QD VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI80_M_u3 VDD net53 QD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI85_M_u2 VDD QD d3 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__icgtp_4 CLK E TE Q VDD VNW VPW VSS
M_MU20 VSS E net50 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU81_M_u2 NCK CLK VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU75_M_u2 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU75_M_u2_22 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU75_M_u2_41 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU75_M_u2_22_37 Q d3 VSS VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU82_M_u3 CK NCK VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MU81_M_u3 VDD CLK NCK VNW pfet_05v0 W=9.2e-07 L=5e-07
M_MI85_M_u1 d3 CLK VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3_3 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3_1 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU75_M_u3_3_28 Q d3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MI82 net50 NCK net53 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI91 net53 CK net033 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI92 net033 QD VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI80_M_u2 VSS net53 QD VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MU82_M_u2 VSS NCK CK VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI85_M_u3 XI85-net6 CLK d3 VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MI85_M_u4 VSS QD XI85-net6 VPW nfet_05v0 W=6.3e-07 L=6e-07
M_MU16 net61 CK net53 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI90 net53 NCK net062 VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI88 net062 QD VDD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI80_M_u3 VDD net53 QD VNW pfet_05v0 W=7.65e-07 L=5e-07
M_MI85_M_u2 VDD QD d3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MU19 net50 TE VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_MI81 VDD TE net58 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_MU17 net58 E net61 VNW pfet_05v0 W=9.25e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
M_i_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VNW VPW VSS
M_i_0_0_x8_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0_x8_1 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0_x8_2 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0_x8_3 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0_x8_4 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0_x8_5 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0_x8_6 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0_x8_7 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0_x8_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_4 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_5 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_6 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0_x8_7 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_12 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_4 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_5 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_6 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_7 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_8 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_9 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_10 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_11 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_16 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_4 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_5 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_6 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_7 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_8 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_9 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_10 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_11 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_12 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_13 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_14 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_15 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_12 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_13 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_14 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_15 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_20 I ZN VDD VNW VPW VSS
M_i_0_0 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_4 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_5 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_6 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_7 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_8 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_9 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_10 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_11 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_12 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_13 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_14 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_15 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_16 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_17 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_18 ZN I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_19 VSS I ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_4 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_5 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_6 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_7 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_8 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_9 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_10 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_11 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_12 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_13 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_14 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_15 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_16 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_17 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_18 ZN I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_19 VDD I ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__invz_1 EN I ZN VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=3.6e-07 L=6e-07
M_mn3 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17 VSS NI NI_N VPW nfet_05v0 W=3.6e-07 L=6e-07
M_Mn_inv NI I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=6.2e-07 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=6.2e-07 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=6.2e-07 L=5e-07
M_mp4 VDD NI_P ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp14 VDD NI NI_P VNW pfet_05v0 W=6.2e-07 L=5e-07
M_Mp_inv NI I VDD VNW pfet_05v0 W=6.2e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__invz_2 EN I ZN VDD VNW VPW VSS
M_XX27 VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX44 NI_N NEN VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX36 NI_P EN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX43 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX22_4 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv NI I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_XX28 VDD EN NEN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_XX45 NI_P EN VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_XX39 NI_N NEN NI_P VNW pfet_05v0 W=1.095e-06 L=5e-07
M_XX46 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_XX21 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_XX21_5 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_Mp_inv NI I VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__invz_3 EN I ZN VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv VSS I NI VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17 NI_N NI VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_mn17_1 VSS NI NI_N VPW nfet_05v0 W=5.4e-07 L=6e-07
M_mn3 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_2 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv VDD I NI VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp14 NI_P NI VDD VNW pfet_05v0 W=1.005e-06 L=5e-07
M_mp14_1 VDD NI NI_P VNW pfet_05v0 W=1.005e-06 L=5e-07
M_mp4 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_1 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_2 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__invz_4 EN I ZN VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv VSS I NI VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17 NI_N NI VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv VDD I NI VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp14 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__invz_8 EN I ZN VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv1 NI I VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_Mn_inv2 VSS I NI VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn17 NI_N NI VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn17_9 VSS NI NI_N VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn17_10 NI_N NI VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn17_9_17 VSS NI NI_N VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn3 ZN NI_N VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn3_1 VSS NI_N ZN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn3_49 ZN NI_N VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn3_1_25 VSS NI_N ZN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn3_99 ZN NI_N VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn3_1_33 VSS NI_N ZN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn3_49_88 ZN NI_N VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mn3_1_25_34 VSS NI_N ZN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv1 NI I VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv2 VDD I NI VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp14 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_11 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10_8 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_58 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_106 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56_111 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57_75 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__invz_12 EN I ZN VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv1 VSS I NI VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv2 NI I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv3 VSS I NI VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17 NI_N NI VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10 NI_N NI VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10_0 NI_N NI VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17_30 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_89 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_34 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_80 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_35 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_99 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_33 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_88 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_34 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv1 VDD I NI VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv2 NI I VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv3 VDD I NI VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp14 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_11 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10_8 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_11_21 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10_8_17 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_57 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_96 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56_105 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57_69 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_58 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_106 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56_111 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57_75 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__invz_16 EN I ZN VDD VNW VPW VSS
M_mn VSS EN NEN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv1 NI I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv2 VSS I NI VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv3 NI I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_Mn_inv4 VSS I NI VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17 NI_N NI VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10 NI_N NI VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_34 NI_N NI VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_41 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_10_30 NI_N NI VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn17_9_17_61 VSS NI NI_N VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_118 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_65 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_181 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_137 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_99_125 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_33_198 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_88_82 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_34_75 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_99 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_33 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_49_88 ZN NI_N VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mn3_1_25_34 VSS NI_N ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_mp VDD EN NEN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp7 NI_P EN VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv1 NI I VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv2 VDD I NI VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv3 NI I VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_Mp_inv4 VDD I NI VNW pfet_05v0 W=1.095e-06 L=5e-07
M_mp14 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_11 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10_8 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_7 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10_32 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_11_55 NI_P NI VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp14_10_8_20 VDD NI NI_P VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_153 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_126 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56_133 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57_97 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_58_95 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_106_111 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56_111_134 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57_75_85 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_58 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_106 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_56_111 ZN NI_P VDD VNW pfet_05v0 W=1.18e-06 L=5e-07
M_mp4_12_57_75 VDD NI_P ZN VNW pfet_05v0 W=1.18e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
M_tn0 VSS E net4 VPW nfet_05v0 W=4.6e-07 L=6e-07
M_tn8 net7 net4 VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn4 VSS D net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net5 net7 net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn1 net2 net4 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn2 net2 net6 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn3 net6 net5 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn6 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp0 VDD E net4 VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp8 net7 net4 VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp5 VDD D net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net1 net4 net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 net5 net7 net0 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 net0 net6 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp3 net6 net5 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp6 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latq_2 D E Q VDD VNW VPW VSS
M_tn0 VSS E net4 VPW nfet_05v0 W=4.6e-07 L=6e-07
M_tn8 net7 net4 VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn4 VSS D net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net5 net7 net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn1 net2 net4 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn2 net2 net6 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn3 net6 net5 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn6_30 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp0 VDD E net4 VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp8 net7 net4 VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp5 VDD D net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net1 net4 net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 net5 net7 net0 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 net0 net6 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp3 net6 net5 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp6_31 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp6 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latq_4 D E Q VDD VNW VPW VSS
M_tn0 VSS E net4 VPW nfet_05v0 W=4.6e-07 L=6e-07
M_tn8 net7 net4 VSS VPW nfet_05v0 W=3.9e-07 L=6e-07
M_tn4 VSS D net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net5 net7 net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn1 net2 net4 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn2 net2 net6 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn3 net6 net5 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn3_94 net6 net5 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn6_30_66 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6_46 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6_30 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn6 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp0 VDD E net4 VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp8 net7 net4 VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp5 VDD D net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net1 net4 net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 net5 net7 net0 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 net0 net6 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp3 net6 net5 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp3_85 net6 net5 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp6_31_68 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp6_71 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp6_31 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp6 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latrnq_1 D E RN Q VDD VNW VPW VSS
M_tn3 net7 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 net1 RN VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn9 net2 D net1 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn8 net2 E net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn7 net3 net7 net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net5 net0 net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn0 VSS RN net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net0 net3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn4 net6 net0 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn1 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net7 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp8 VDD RN net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net8 D VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net3 net7 net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net9 E net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net9 net0 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net0 net3 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7 net6 net0 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp0 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latrnq_2 D E RN Q VDD VNW VPW VSS
M_tn3 net7 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 net1 RN VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn9 net2 D net1 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn8 net2 E net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn7 net3 net7 net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net5 net0 net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn0 VSS RN net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net0 net3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn4 net6 net0 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn1 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1_38 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net7 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp8 VDD RN net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net8 D VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net3 net7 net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net9 E net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net9 net0 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net0 net3 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7 net6 net0 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp0 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_27 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latrnq_4 D E RN Q VDD VNW VPW VSS
M_tn3 net7 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 net1 RN VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn9 net2 D net1 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn8 net2 E net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn7 net3 net7 net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net5 net0 net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn0 VSS RN net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net0 net3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn6_109 net0 net3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn4 net6 net0 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn4_77 net6 net0 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn1 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1_38 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1_15 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1_38_14 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net7 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp8 VDD RN net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net8 D VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net3 net7 net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net9 E net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net9 net0 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net0 net3 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp9_110 net0 net3 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7 net6 net0 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7_78 net6 net0 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp0 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_27 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_24 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_27_20 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latrsnq_1 D E RN SETN Q VDD VNW VPW VSS
M_tn3 net8 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn9 net2 RN VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn8 net3 D net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn7 net3 E net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net4 net8 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net6 net1 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn0 VSS RN net6 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn11 VSS net4 net0 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 net0 SETN net1 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn4 net7 net1 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn1 Q net7 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net8 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp8 VDD RN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net9 D VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net4 net8 net9 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net10 E net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net10 net1 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 VDD net4 net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net1 SETN VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7 net7 net1 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp0 Q net7 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latrsnq_2 D E RN SETN Q VDD VNW VPW VSS
M_tn3 net8 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn9 net2 RN VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn8 net3 D net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn7 net3 E net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net4 net8 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net6 net1 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn0 VSS RN net6 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn11 VSS net4 net0 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 net0 SETN net1 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn4 net7 net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1 Q net7 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1_19 Q net7 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net8 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp8 VDD RN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net9 D VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net4 net8 net9 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net10 E net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net10 net1 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 VDD net4 net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net1 SETN VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7 net7 net1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0 Q net7 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_9 Q net7 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latrsnq_4 D E RN SETN Q VDD VNW VPW VSS
M_tn3 net8 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn9 net2 RN VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn8 net3 D net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn7 net3 E net4 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net4 net8 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net6 net1 net5 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn0 VSS RN net6 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn11 VSS net4 net0 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn10 net0 SETN net1 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn4_44 net7 net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn4 net7 net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1 Q net7 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1_19 Q net7 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1_18 Q net7 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn1_19_0 Q net7 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net8 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp8 VDD RN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net9 D VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net4 net8 net9 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net10 E net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net10 net1 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 VDD net4 net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net1 SETN VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7_47 net7 net1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp7 net7 net1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0 Q net7 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_9 Q net7 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_26 Q net7 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_9_34 Q net7 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latsnq_1 D E SETN Q VDD VNW VPW VSS
M_tn2 net6 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn7 VSS D net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net3 E net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net4 net6 net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn4 net4 net1 VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn9 VSS net3 net0 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn8 net0 SETN net1 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn3 net5 net1 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn0 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net6 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp6 VDD D net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net7 net6 net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net3 E net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net8 net1 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 VDD net3 net1 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp8 net1 SETN VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7 net5 net1 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp0 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latsnq_2 D E SETN Q VDD VNW VPW VSS
M_tn2 net6 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn7 VSS D net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net3 E net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net4 net6 net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn4 net4 net1 VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn9 VSS net3 net0 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn8 net0 SETN net1 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn3 net5 net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn0 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn0_11 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net6 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp6 VDD D net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net7 net6 net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net3 E net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net8 net1 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 VDD net3 net1 VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp8 net1 SETN VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp7 net5 net1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_8 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__latsnq_4 D E SETN Q VDD VNW VPW VSS
M_tn2 net6 E VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn7 VSS D net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn6 net3 E net2 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn5 net4 net6 net3 VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn4 net4 net1 VSS VPW nfet_05v0 W=3.95e-07 L=6e-07
M_tn9 VSS net3 net0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn8 net0 SETN net1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn3_56 net5 net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn3 net5 net1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn0 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn0_11 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn0_12 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn0_11_1 Q net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp2 net6 E VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp6 VDD D net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net7 net6 net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 net3 E net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net8 net1 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 VDD net3 net1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp8 net1 SETN VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp7_53 net5 net1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp7 net5 net1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_8 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_32 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp0_8_30 Q net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__mux2_1 I0 I1 S Z VDD VNW VPW VSS
M_MN2 VSS int04 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN4 net_1 I1 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_MN8 int04 S net_1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_MN7 net_3 sel1_n int04 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_MN3 VSS I0 net_3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_MN1 sel1_n S VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_MP5 VDD int04 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP4 net_0 I1 VDD VNW pfet_05v0 W=6.15e-07 L=5e-07
M_MP8 int04 sel1_n net_0 VNW pfet_05v0 W=6.15e-07 L=5e-07
M_MP7 net_2 S int04 VNW pfet_05v0 W=6.15e-07 L=5e-07
M_MP3 VDD I0 net_2 VNW pfet_05v0 W=6.15e-07 L=5e-07
M_MP1 sel1_n S VDD VNW pfet_05v0 W=6.15e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
M_MN2_12 VSS int04 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN2 VSS int04 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN4 net_1 I1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN8 int04 S net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN7 net_3 sel1_n int04 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN3 VSS I0 net_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN1 sel1_n S VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MP5_6 VDD int04 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP5 VDD int04 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP4 net_0 I1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP8 int04 sel1_n net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP7 net_2 S int04 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP3 VDD I0 net_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP1 sel1_n S VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
M_MN2_12_7 VSS int04 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN2_8 VSS int04 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN2_12 VSS int04 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN2 VSS int04 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN4 net_1 I1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN8 int04 S net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN7 net_3 sel1_n int04 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN3 VSS I0 net_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MN1 sel1_n S VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_MP5_6_5 VDD int04 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP5_0 VDD int04 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP5_6 VDD int04 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP5 VDD int04 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP4 net_0 I1 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP8 int04 sel1_n net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP7 net_2 S int04 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP3 VDD I0 net_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_MP1 sel1_n S VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
M_MN5 int01 I2 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN9 int02 sel1_n int01 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN10 int07 S0 int02 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN6 VSS I3 int07 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_instance_22 Z int03 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN12 int03 S1 int02 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN11 int04 sel2_n int03 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN2 VSS S1 sel2_n VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN4 int06 I1 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN8 int04 S0 int06 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN7 int05 sel1_n int04 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN3 VSS I0 int05 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN1 sel1_n S0 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MP2 int01 I2 VDD VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP9 int02 S0 int01 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP10 int07 sel1_n int02 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP6 VDD I3 int07 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_instance_1 Z int03 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP12 int03 sel2_n int02 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP11 int04 S1 int03 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP5 VDD S1 sel2_n VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP4 int06 I1 VDD VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP8 int04 sel1_n int06 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP7 int05 S0 int04 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP3 VDD I0 int05 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_MP1 sel1_n S0 VDD VNW pfet_05v0 W=5.65e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
M_MN5 int01 I2 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN9 int02 sel1_n int01 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN10 int07 S0 int02 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN6 VSS I3 int07 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_instance_22 Z int03 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_instance_22_11 Z int03 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN12 int03 S1 int02 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN11 int04 sel2_n int03 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN2 VSS S1 sel2_n VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN4 int06 I1 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN8 int04 S0 int06 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN7 int05 sel1_n int04 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN3 VSS I0 int05 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN1 sel1_n S0 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MP2 int01 I2 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP9 int02 S0 int01 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP10 int07 sel1_n int02 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP6 VDD I3 int07 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_instance_1 Z int03 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_instance_1_6 Z int03 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP12 int03 sel2_n int02 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP11 int04 S1 int03 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP5 VDD S1 sel2_n VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP4 int06 I1 VDD VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP8 int04 sel1_n int06 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP7 int05 S0 int04 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP3 VDD I0 int05 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP1 sel1_n S0 VDD VNW pfet_05v0 W=5.95e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
M_MN5 int01 I2 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN9 int02 sel1_n int01 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN10 int07 S0 int02 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN6 VSS I3 int07 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_instance_22 Z int03 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_instance_22_11 Z int03 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_instance_22_18 Z int03 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_instance_22_11_19 Z int03 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_MN12 int03 S1 int02 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN11 int04 sel2_n int03 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN2 VSS S1 sel2_n VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN4 int06 I1 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN8 int04 S0 int06 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN7 int05 sel1_n int04 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN3 VSS I0 int05 VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MN1 sel1_n S0 VSS VPW nfet_05v0 W=3.65e-07 L=6e-07
M_MP2 int01 I2 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP9 int02 S0 int01 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP10 int07 sel1_n int02 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP6 VDD I3 int07 VNW pfet_05v0 W=7.8e-07 L=5e-07
M_instance_1 Z int03 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_instance_1_6 Z int03 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_instance_1_9 Z int03 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_instance_1_6_3 Z int03 VDD VNW pfet_05v0 W=7.8e-07 L=5e-07
M_MP12 int03 sel2_n int02 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP11 int04 S1 int03 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP5 VDD S1 sel2_n VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP4 int06 I1 VDD VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP8 int04 sel1_n int06 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP7 int05 S0 int04 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP3 VDD I0 int05 VNW pfet_05v0 W=5.95e-07 L=5e-07
M_MP1 sel1_n S0 VDD VNW pfet_05v0 W=5.95e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
M_i_1 net_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 ZN A2 VDD VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_2 VDD A1 ZN VNW pfet_05v0 W=1.13e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
M_i_1_1 net_0_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0_1 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 VSS A2 net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 ZN A2 VDD VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_2_1 VDD A1 ZN VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_2_0 ZN A1 VDD VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_3_0 VDD A2 ZN VNW pfet_05v0 W=1.13e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
M_i_1_3 net_0_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 ZN A1 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 net_0_1 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 VSS A2 net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0_2 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0_3 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 VSS A2 net_0_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_3 ZN A2 VDD VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_2_3 VDD A1 ZN VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_2_2 ZN A1 VDD VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_3_2 VDD A2 ZN VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_3_1 ZN A2 VDD VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_2_1 VDD A1 ZN VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_2_0 ZN A1 VDD VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_3_0 VDD A2 ZN VNW pfet_05v0 W=1.13e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_2 net_1 A3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 net_0 A2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5 ZN A3 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_4 VDD A2 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_3 ZN A1 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_2_1 net_1_0 A3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0_0 A2 net_1_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0_1 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_1_1 A2 net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 VSS A3 net_1_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 ZN A3 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_4_0 VDD A2 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_3_0 ZN A1 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_3_1 VDD A1 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_4_1 ZN A2 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_5_0 VDD A3 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_1_3 net_1_3 A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 VSS A3 net_1_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_1_2 A3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_0 A2 net_1_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_1_1 A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 VSS A3 net_1_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 net_1_0 A3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0_0 A2 net_1_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 ZN A1 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_3 ZN A2 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_5_0 VDD A3 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_5_1 ZN A3 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_4_2 VDD A2 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_4_1 ZN A2 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_5_2 VDD A3 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_5_3 ZN A3 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_4_0 VDD A2 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_3_3 ZN A1 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_3_2 VDD A1 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_3_1 ZN A1 VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_3_0 VDD A1 ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
M_i_3 net_2 A4 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_1 A3 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 net_0 A2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7 ZN A4 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_6 VDD A3 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_5 ZN A2 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_4 VDD A1 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
M_i_3_0 net_2_0 A4 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_1_0 A3 net_2_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0_0 A2 net_1_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0_1 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_1_1 A2 net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_2_1 A3 net_1_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 VSS A4 net_2_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7_0 VDD A4 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_6_0 ZN A3 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_5_0 VDD A2 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_4_0 ZN A1 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_4_1 VDD A1 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_5_1 ZN A2 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_6_1 VDD A3 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_7_1 ZN A4 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
M_i_2_3 net_2_3 A3 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_3 VSS A4 net_2_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 net_2_2 A4 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_1 A3 net_2_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_2_1 A3 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 VSS A4 net_2_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_2_0 A4 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_1_0 A3 net_2_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 net_0_3 A2 net_1_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 ZN A1 net_0_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 net_0_2 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_1 A2 net_0_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0_1 A2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_1 A2 net_0_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_3 ZN A3 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_7_3 VDD A4 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_7_2 ZN A4 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_6_2 VDD A3 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_6_1 ZN A3 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_7_1 VDD A4 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_7_0 ZN A4 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_6_0 VDD A3 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_5_3 ZN A2 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_4_3 VDD A1 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_4_2 ZN A1 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_5_2 VDD A2 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_5_1 ZN A2 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_4_1 VDD A1 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_4_0 ZN A1 VDD VNW pfet_05v0 W=8.45e-07 L=5e-07
M_i_5_0 VDD A2 ZN VNW pfet_05v0 W=8.45e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
M_i_1 ZN A2 VSS VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_0 VSS A1 ZN VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_3 net_0 A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_2 ZN A1 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
M_i_1_1 ZN A2 VSS VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_0_1 VSS A1 ZN VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_0_0 ZN A1 VSS VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_1_0 VSS A2 ZN VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_3_1 net_0_0 A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_2_1 ZN A1 net_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_2_0 net_0_1 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0 VDD A2 net_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
M_i_1_3 ZN A2 VSS VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_0_3 VSS A1 ZN VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_0_2 ZN A1 VSS VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_1_2 VSS A2 ZN VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_1_1 ZN A2 VSS VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_0_1 VSS A1 ZN VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_0_0 ZN A1 VSS VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_1_0 VSS A2 ZN VPW nfet_05v0 W=5.65e-07 L=6e-07
M_i_3_3 net_0_0 A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_2_3 ZN A1 net_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_2_2 net_0_1 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_2 VDD A2 net_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_1 net_0_2 A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_2_1 ZN A1 net_0_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_2_0 net_0_3 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0 VDD A2 net_0_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_2 ZN A3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_1 VSS A2 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0 ZN A1 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_5 net_1 A3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4 net_0 A2 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3 ZN A1 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_2_1 VSS A3 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_1_0 ZN A2 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0_0 VSS A1 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0_1 ZN A1 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_1_1 VSS A2 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_2_0 ZN A3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_5_1 net_1_0 A3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_0 net_0_0 A2 net_1_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0 ZN A1 net_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_1 net_0_1 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_1 net_1_1 A2 net_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_0 VDD A3 net_1_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_1_3 ZN A2 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_2_0 VSS A3 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_2_1 ZN A3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_1_2 VSS A2 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_1_1 ZN A2 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_2_2 VSS A3 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_2_3 ZN A3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_1_0 VSS A2 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0_3 ZN A1 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0_2 VSS A1 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0_1 ZN A1 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0_0 VSS A1 ZN VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_4_3 net_1_3 A2 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_0 VDD A3 net_1_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_1 net_1_2 A3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_2 net_0 A2 net_1_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_1 net_1_1 A2 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_2 VDD A3 net_1_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_3 net_1_0 A3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_0 net_0_0 A2 net_1_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_3 ZN A1 net_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_2 net_0 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_1 ZN A1 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3_0 net_0 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
M_i_3 ZN A4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 VSS A3 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1 ZN A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 VSS A1 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_7 net_2 A4 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6 net_1 A3 net_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5 net_0 A2 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4 ZN A1 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
M_i_2_1 ZN A3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_1 VSS A4 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_0 ZN A4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0 VSS A3 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1_1 ZN A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_1 VSS A1 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_0 ZN A1 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1_0 VSS A2 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_6_1 net_2_1 A3 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 VDD A4 net_2_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 net_2_0 A4 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0 net_1_0 A3 net_2_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_1 net_0_1 A2 net_1_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_1 ZN A1 net_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_0 net_0_0 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_0 net_1 A2 net_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
M_i_2_3 ZN A3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_3 VSS A4 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_2 ZN A4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_2 VSS A3 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_1 ZN A3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_1 VSS A4 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3_0 ZN A4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2_0 VSS A3 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1_3 ZN A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_3 VSS A1 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_2 ZN A1 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1_2 VSS A2 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1_1 ZN A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_1 VSS A1 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0_0 ZN A1 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1_0 VSS A2 ZN VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_6_3 net_2_3 A3 net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7_3 VDD A4 net_2_3 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7_2 net_2_2 A4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_2 net_1 A3 net_2_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_1 net_2_1 A3 net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7_1 VDD A4 net_2_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_7_0 net_2_0 A4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_6_0 net_1_0 A3 net_2_0 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_3 net_0_3 A2 net_1_0 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4_3 ZN A1 net_0_3 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4_2 net_0_2 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_2 net_1 A2 net_0_2 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_1 net_0_1 A2 net_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4_1 ZN A1 net_0_1 VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_4_0 net_0_0 A1 ZN VNW pfet_05v0 W=1.215e-06 L=5e-07
M_i_5_0 net_1 A2 net_0_0 VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
M_i_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 VSS B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4 net_1 A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3 ZN A1 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5 VDD B ZN VNW pfet_05v0 W=1.13e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
M_i_2_1 VSS B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 B VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 ZN B VDD VNW pfet_05v0 W=9.55e-07 L=5e-07
M_i_5_0 VDD B ZN VNW pfet_05v0 W=9.55e-07 L=5e-07
M_i_4_1 net_1_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3_1 ZN A1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3_0 net_1_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 VDD A2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
M_i_1_3 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 VSS B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_0 B VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 B VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_3 net_1_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3_3 ZN A1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3_2 net_1_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_2 VDD A2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_1 net_1_2 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3_1 ZN A1 net_1_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3_0 net_1_3 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 VDD A2 net_1_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_3 ZN B VDD VNW pfet_05v0 W=9.55e-07 L=5e-07
M_i_5_2 VDD B ZN VNW pfet_05v0 W=9.55e-07 L=5e-07
M_i_5_1 ZN B VDD VNW pfet_05v0 W=9.55e-07 L=5e-07
M_i_5_0 VDD B ZN VNW pfet_05v0 W=9.55e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
M_i_3 VSS B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_0 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7 net_2 B2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6 ZN B1 net_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4 net_1 A1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5 VDD A2 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
M_i_3_1 VSS B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_0 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 VSS B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_0 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7_1 net_2_0 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 ZN B1 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_2_1 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 VDD B2 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 net_1_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_1 ZN A1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 net_1_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 VDD A2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
M_i_3_3 VSS B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 net_0 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 VSS B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 net_0 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 VSS B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_0 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 VSS B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_0 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7_3 net_2_0 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_3 ZN B1 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_2 net_2_1 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_2 VDD B2 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 net_2_2 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 ZN B1 net_2_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_2_3 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 VDD B2 net_2_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 net_1_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 ZN A1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_1 net_1_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 VDD A2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_2 net_1_2 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_2 ZN A1 net_1_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_3 net_1_3 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_3 VDD A2 net_1_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
M_i_3 net_0 B VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_1 net_0 A2 ZN VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_2 ZN A3 net_0 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_i_7 ZN B VDD VNW pfet_05v0 W=1.13e-06 L=5e-07
M_i_4 net_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5 net_2 A2 net_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6 VDD A3 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
M_i_3_1 VSS B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_0 B VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 ZN A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 A3 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7_1 ZN B VDD VNW pfet_05v0 W=1.08e-06 L=5e-07
M_i_7_0 VDD B ZN VNW pfet_05v0 W=1.08e-06 L=5e-07
M_i_6_1 net_2_0 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 net_1_0 A2 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_1 ZN A1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 net_1_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 net_2_1 A2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 VDD A3 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
M_i_2_3 ZN A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_0 A3 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 ZN A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 A3 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_3 VSS B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 net_0 B VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 VSS B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_0 B VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_3 VDD A3 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_2 net_2 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 VDD A3 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_2_0 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_3 net_1_0 A2 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_3 ZN A1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_2 net_1_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_2 net_2 A2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 net_1_2 A2 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_1 ZN A1 net_1_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 net_1_3 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 net_2 A2 net_1_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_3 ZN B VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_2 VDD B ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 ZN B VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 VDD B ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
M_i_4 net_0 A3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VSS A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_0 A1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 net_0 B2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9 net_3 A3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8 net_2 A2 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7 ZN A1 net_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5 net_1 B1 ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6 VDD B2 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
M_i_4_1 VSS A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 A1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 net_0 A3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0 B2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9_1 net_3_0 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_1 net_2_0 A2 net_3_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 ZN A1 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 net_2_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_0 net_3_1 A2 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_0 VDD A3 net_3_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_1_0 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 ZN B1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 net_1_1 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 VDD B2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
M_i_3_3 VSS A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_3 net_0 A3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_2 VSS A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 net_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 VSS A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_1 net_0 A3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 VSS A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_0 A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 VSS A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_0 A1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 A1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 ZN B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 net_0 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_0 B2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 B1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 B2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8_3 net_3_0 A2 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_3 VDD A3 net_3_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_2 net_3_1 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_2 net_2 A2 net_3_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_1 net_3_2 A2 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_1 VDD A3 net_3_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_0 net_3_3 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_0 net_2_0 A2 net_3_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_3 ZN A1 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_2 net_2 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 ZN A1 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 net_2 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_3 net_1_0 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_3 ZN B1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_2 net_1_1 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_2 VDD B2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 net_1_2 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 ZN B1 net_1_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 net_1_3 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 VDD B2 net_1_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
M_i_5 net_0 B3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4 VSS B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 net_0 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 ZN A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_11 net_4 B3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10 net_3 B2 net_4 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9 ZN B1 net_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6 net_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7 net_2 A2 net_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8 VDD A3 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai33_2 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
M_i_5_0 VSS B3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_1 net_0 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 VSS B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_0 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 VSS B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 net_0 B3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 ZN A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_0 A3 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_11_0 net_4_0 B3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_1 net_3_0 B2 net_4_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_1 ZN B1 net_3_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_0 net_3_1 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_0 net_4_1 B2 net_3_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_1 VDD B3 net_4_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_0 net_2_0 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 net_1_0 A2 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 ZN A1 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_1_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 net_2_1 A2 net_1_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_1 VDD A3 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
M_i_4_0 VSS B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_0 net_0 B3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 VSS B3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_1 net_0 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_2 VSS B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_2 net_0 B3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_3 VSS B3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_3 net_0 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_0 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 VSS B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_3 net_0 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 net_0 A3 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 ZN A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_0 A3 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 ZN A3 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10_0 net_4_0 B2 net_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_0 VDD B3 net_4_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_1 net_4_1 B3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_1 net_3 B2 net_4_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_2 net_4_2 B2 net_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_2 VDD B3 net_4_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_3 net_4_3 B3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_3 net_3_0 B2 net_4_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_0 ZN B1 net_3_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_1 net_3 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_2 ZN B1 net_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_3 net_3 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 ZN A1 net_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 net_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_2 ZN A1 net_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_3 net_1_0 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_3 net_2_0 A2 net_1_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_3 VDD A3 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_2 net_2_1 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_2 net_1 A2 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 net_2_2 A2 net_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_1 VDD A3 net_2_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_0 net_2_3 A3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 net_1 A2 net_2_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
M_i_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_1 B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VSS C net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5 net_2 A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4 ZN A1 net_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6 VDD B ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_7 ZN C VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_1_0 B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS C net_1_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_1_1 C VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_0 B net_1_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 net_2_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_1 ZN A1 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 net_2_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 VDD A2 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 ZN B VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_7_0 VDD C ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_7_1 ZN C VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_6_1 VDD B ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
M_i_1_3 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_1_0 B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS C net_1_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_1_1 C VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_0 B net_1_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_1_2 B net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 VSS C net_1_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_3 net_1_3 C VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 net_0 B net_1_3 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_3 net_2_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_3 ZN A1 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_2 net_2_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_2 VDD A2 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 net_2_2 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_1 ZN A1 net_2_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4_0 net_2_3 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 VDD A2 net_2_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 ZN B VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_7_0 VDD C ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_7_1 ZN C VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_6_1 VDD B ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_6_2 ZN B VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_7_2 VDD C ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_7_3 ZN C VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_6_3 VDD B ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
M_i_4 VSS B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 net_1 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_0 C net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9 net_3 B2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8 ZN B1 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7 VDD C ZN VNW pfet_05v0 W=9.45e-07 L=5e-07
M_i_6 net_2 A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5 ZN A1 net_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
M_i_2_1 net_1 C net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_1 VSS B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_1 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS B1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 net_1 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 C net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7_1 VDD C ZN VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_9_1 net_3_0 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_1 ZN B1 net_3_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_0 net_3_1 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_0 VDD B2 net_3_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 ZN C VDD VNW pfet_05v0 W=9.85e-07 L=5e-07
M_i_5_1 net_2_0 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 VDD A2 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_2_1 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 ZN A1 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
M_i_3_3 net_1 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_3 VSS B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_2 net_1 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 VSS B1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_1 B1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_1 VSS B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 net_1 B2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS B1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 net_1 C net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_0 C net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_1 C net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_0 C net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8_3 net_3_0 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_3 VDD B2 net_3_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_2 net_3_1 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_2 ZN B1 net_3_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_1 net_3_2 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_1 VDD B2 net_3_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_0 net_3_3 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_0 ZN B1 net_3_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_3 VDD C ZN VNW pfet_05v0 W=9.35e-07 L=5e-07
M_i_7_2 ZN C VDD VNW pfet_05v0 W=9.35e-07 L=5e-07
M_i_7_1 VDD C ZN VNW pfet_05v0 W=9.35e-07 L=5e-07
M_i_7_0 ZN C VDD VNW pfet_05v0 W=9.35e-07 L=5e-07
M_i_5_3 net_2_0 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_3 VDD A2 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_2 net_2_1 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_2 ZN A1 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_1 net_2_2 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 VDD A2 net_2_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_2_3 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5_0 ZN A1 net_2_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
M_i_5 net_1 C2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4 VSS C1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_1 B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 net_0 B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_11 net_4 C2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10 ZN C1 net_4 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8 net_3 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9 VDD B2 net_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7 net_2 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6 ZN A1 net_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
M_i_4_1 net_1 C1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 VSS C2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_0 net_1 C2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 VSS C1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_1 B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_0 B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_1 B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_0 B1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10_1 net_4_1 C1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_1 VDD C2 net_4_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_0 net_4_0 C2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_0 ZN C1 net_4_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_0 net_3_1 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_0 VDD B2 net_3_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_1 net_3_0 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_1 ZN B1 net_3_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_2_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 VDD A2 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 net_2_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 ZN A1 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
M_i_4_3 net_1 C1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_3 VSS C2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_2 net_1 C2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_2 VSS C1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_1 net_1 C1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 VSS C2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_0 net_1 C2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4_0 VSS C1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 net_1 B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 net_0 B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_1 net_1 B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 net_0 B1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_2 net_1 B1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_2 net_0 B2 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_3 net_1 B2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_3 net_0 B1 net_1 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_2 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1_3 ZN A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 net_0 A1 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10_3 net_4_3 C1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_3 VDD C2 net_4_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_2 net_4_2 C2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_2 ZN C1 net_4_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_1 net_4_1 C1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_1 VDD C2 net_4_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11_0 net_4_0 C2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10_0 ZN C1 net_4_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_0 net_3_3 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_0 VDD B2 net_3_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_1 net_3_2 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_1 ZN B1 net_3_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_2 net_3_1 B1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_2 VDD B2 net_3_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9_3 net_3_0 B2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_8_3 ZN B1 net_3_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_0 net_2_3 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_0 VDD A2 net_2_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 net_2_2 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_1 ZN A1 net_2_2 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_2 net_2_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_2 VDD A2 net_2_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_3 net_2_0 A2 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6_3 ZN A1 net_2_0 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
M_i_2 Z_neg A1 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 VSS A2 Z_neg VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4 net_0 A1 Z_neg VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_5 VDD A2 net_0 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
M_i_2 Z_neg A1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VSS A2 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_4 net_0 A1 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5 VDD A2 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
M_i_3_1 Z_neg A2 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_1 VSS A1 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2_0 Z_neg A1 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3_0 VSS A2 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5_1 net_0_1 A2 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_1 Z_neg A1 net_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4_0 net_0_0 A1 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_0 VDD A2 net_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
M_i_2 VSS A1 Z_neg VPW nfet_05v0 W=4e-07 L=6e-07
M_i_3 Z_neg A2 VSS VPW nfet_05v0 W=4e-07 L=6e-07
M_i_4 VSS A3 Z_neg VPW nfet_05v0 W=4e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5 net_0 A1 Z_neg VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_6 net_1 A2 net_0 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_7 VDD A3 net_1 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
M_i_2 VSS A1 Z_neg VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_3 Z_neg A2 VSS VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_4 VSS A3 Z_neg VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_5 net_0 A1 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6 net_1 A2 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7 VDD A3 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
M_i_4_0 Z_neg A3 VSS VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_3_1 VSS A2 Z_neg VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_2_1 Z_neg A1 VSS VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_2_0 VSS A1 Z_neg VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_3_0 Z_neg A2 VSS VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_4_1 VSS A3 Z_neg VPW nfet_05v0 W=6.65e-07 L=6e-07
M_i_0_3 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7_0 net_1_1 A3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_1 net_0_1 A2 net_1_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_1 Z_neg A1 net_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5_0 net_0_0 A1 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0 net_1_0 A2 net_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 VDD A3 net_1_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
M_i_2 Z_neg A1 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_3 VSS A2 Z_neg VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_4 Z_neg A3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_5 VSS A4 Z_neg VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6 net_0 A1 Z_neg VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_7 net_1 A2 net_0 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_8 net_2 A3 net_1 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_9 VDD A4 net_2 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
M_i_2 Z_neg A1 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_3 VSS A2 Z_neg VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_4 Z_neg A3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_5 VSS A4 Z_neg VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6 net_0 A1 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7 net_1 A2 net_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8 net_2 A3 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9 VDD A4 net_2 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
M_i_5_1_x2_1 Z_neg A4 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_4_1_x2_1 VSS A3 Z_neg VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_3_1_x2_1 Z_neg A2 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_2_1_x2_1 VSS A1 Z_neg VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_2_1_x2_0 Z_neg A1 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_3_1_x2_0 VSS A2 Z_neg VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_4_1_x2_0 Z_neg A3 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_5_1_x2_0 VSS A4 Z_neg VPW nfet_05v0 W=4.65e-07 L=6e-07
M_i_0_3_x4_3 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3_x4_2 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3_x4_1 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3_x4_0 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9_0_m2_1 net_2_0_1 A4 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8_0_m2_1 net_1_0_1 A3 net_2_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0_m2_1 net_0_0_1 A2 net_1_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0_m2_1 Z_neg A1 net_0_0_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6_0_m2_0 net_0_0_0 A1 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0_m2_0 net_1_0_0 A2 net_0_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_8_0_m2_0 net_2_0_0 A3 net_1_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9_0_m2_0 VDD A4 net_2_0_0 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3_x4_3 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3_x4_2 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3_x4_1 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3_x4_0 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffq_1 D SE SI CLK Q VDD VNW VPW VSS
M_tn14 net8 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net12 SI VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net12 SE net6 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net6 net8 net9n VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 VSS D net9n VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn9 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn11 net6 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net5 cki net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 VSS net10 net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 net5 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 cki net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net7 ncki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 VSS net1 net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net1 net0 VSS VPW nfet_05v0 W=4.35e-07 L=6e-07
M_tn6 Q net1 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp14 net8 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net3 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp12 net2 net8 net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 net9p SE net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 VDD D net9p VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 ncki CLK VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp9 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp11 net5 cki net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp0 net4 ncki net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 VDD net10 net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp15 net10 net5 VDD VNW pfet_05v0 W=6.3e-07 L=5.1e-07
M_tp7 net0 ncki net10 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net7_p cki net0 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 VDD net1 net7_p VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net1 net0 VDD VNW pfet_05v0 W=7.05e-07 L=5e-07
M_tp4 Q net1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffq_2 D SE SI CLK Q VDD VNW VPW VSS
M_tn14 net8 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net12 SI VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net12 SE net6 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net6 net8 net9n VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 VSS D net9n VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn9 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn11 net6 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net5 cki net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 VSS net10 net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 net5 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 cki net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net7 ncki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 VSS net1 net7 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn5 net1 net0 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn6_6 Q net1 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn6 Q net1 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp14 net8 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net3 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp12 net2 net8 net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 net9p SE net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 VDD D net9p VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 ncki CLK VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp9 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp11 net5 cki net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp0 net4 ncki net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 VDD net10 net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp15 net10 net5 VDD VNW pfet_05v0 W=6.3e-07 L=5.1e-07
M_tp7 net0 ncki net10 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net7_p cki net0 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 VDD net1 net7_p VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp3 net1 net0 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp4_12 Q net1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp4 Q net1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffq_4 D SE SI CLK Q VDD VNW VPW VSS
M_tn14 net8 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net12 SI VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net12 SE net6 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net6 net8 net9n VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 VSS D net9n VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn9 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn11 net6 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net5 cki net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 VSS net10 net11 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net10 net5 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 cki net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net7 ncki net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 VSS net1 net7 VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn5 net1 net0 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn6_6_25 Q net1 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn6_5 Q net1 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn6_6 Q net1 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn6 Q net1 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp14 net8 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net3 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp12 net2 net8 net3 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 net9p SE net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 VDD D net9p VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 ncki CLK VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp9 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp11 net5 cki net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp0 net4 ncki net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 VDD net10 net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp15 net10 net5 VDD VNW pfet_05v0 W=6.3e-07 L=5.1e-07
M_tp7 net0 ncki net10 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 net7_p cki net0 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 VDD net1 net7_p VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp3 net1 net0 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp4_12_24 Q net1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp4_16 Q net1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp4_12 Q net1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp4 Q net1 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1 D RN SE SI CLK Q VDD VNW VPW VSS
M_tn17 net3 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS SI net13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net13 SE net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net10 D net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 net5 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn13 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn15 net10 ncki net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 cki net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net8 cki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net11 ncki net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tp17 net3 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 net7 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net6 net3 net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net14 D net6 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp14 VDD SE net14 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp11 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp15 net1 cki net6 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp7 net9 ncki net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 net2 ncki net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net8 cki net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2 D RN SE SI CLK Q VDD VNW VPW VSS
M_tn17 net3 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS SI net13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net13 SE net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net10 D net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 net5 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn13 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn15 net10 ncki net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 cki net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net8 cki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net11 ncki net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn3_17 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tp17 net3 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 net7 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net6 net3 net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net14 D net6 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp14 VDD SE net14 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp11 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp15 net1 cki net6 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp7 net9 ncki net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 net2 ncki net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net8 cki net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp1_16 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4 D RN SE SI CLK Q VDD VNW VPW VSS
M_tn17 net3 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS SI net13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net13 SE net10 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net10 D net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 net5 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn13 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn15 net10 ncki net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 cki net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net12 net2 net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS RN net12 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 VSS net1 net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net8 cki net2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net11 ncki net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net11 net4 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net0 RN VSS VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn4 net4 net8 net0 VPW nfet_05v0 W=5.4e-07 L=6e-07
M_tn3_17_4 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tn3_27 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tn3_17 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tn3 Q net4 VSS VPW nfet_05v0 W=8.1e-07 L=6e-07
M_tp17 net3 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 net7 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net6 net3 net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 net14 D net6 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp14 VDD SE net14 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp11 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp15 net1 cki net6 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp7 net9 ncki net1 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp6 VDD net2 net9 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp12 net9 RN VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp18 VDD net1 net2 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp2 net2 ncki net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp3 net8 cki net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 net11 net4 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp5 net4 RN VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp4 VDD net8 net4 VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp1_16_17 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1_25 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1_16 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
M_tp1 Q net4 VDD VNW pfet_05v0 W=1.215e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1 D RN SE SETN SI CLK Q VDD VNW VPW VSS
M_tn12 net9 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS SI net17 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 net17 SE net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net14 D net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net8 net9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn2 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn8 net14 ncki net3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net3 cki net16 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp12 net9 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp11 net12 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 net10 net9 net12 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp0 net11 D net10 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 VDD SE net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp2 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp10 net3 cki net10 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp7 net13 ncki net3 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp20 net4 ncki net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp19 net5 cki net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=9.2e-07 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2 D RN SE SETN SI CLK Q VDD VNW VPW VSS
M_tn12 net9 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS SI net17 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 net17 SE net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net14 D net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net8 net9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn2 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn8 net14 ncki net3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net3 cki net16 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn19_14 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp12 net9 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp11 net12 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 net10 net9 net12 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp0 net11 D net10 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 VDD SE net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp2 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp10 net3 cki net10 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp7 net13 ncki net3 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp20 net4 ncki net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp19 net5 cki net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp17_7 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4 D RN SE SETN SI CLK Q VDD VNW VPW VSS
M_tn12 net9 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 VSS SI net17 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 net17 SE net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn0 net14 D net8 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn11 net8 net9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn2 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn8 net14 ncki net3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 net3 cki net16 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn6 net15 net4 net16 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS RN net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 net1 SETN net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn16 VSS net6 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 net2 RN VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn17 net6 net5 net2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn19 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn19_14 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn19_12 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn19_14_0 Q net6 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp12 net9 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp11 net12 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 net10 net9 net12 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp0 net11 D net10 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp9 VDD SE net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp2 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp10 net3 cki net10 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp7 net13 ncki net3 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp5 VDD net4 net13 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp6 net13 RN VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp4 VDD net3 net4 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp3 VDD SETN net4 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp20 net4 ncki net5 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp19 net5 cki net7 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp13 net7 SETN VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp14 net7 net6 VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp16 net6 RN VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp15 VDD net5 net6 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp17 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp17_7 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp17_8 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp17_7_4 Q net6 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1 D SE SETN SI CLK Q VDD VNW VPW VSS
M_tn11 net9 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS SI net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 net15 SE net13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 net13 D net16 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net16 net9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn0 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn6 net13 ncki net3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net3 cki net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp11 net9 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 net11 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 net8 net9 net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 net12 D net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp7 VDD SE net12 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp0 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp9 net3 cki net8 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp6 net10 ncki net3 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp18 net5 ncki net4 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp17 net7 cki net5 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2 D SE SETN SI CLK Q VDD VNW VPW VSS
M_tn11 net9 SE VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn7 VSS SI net15 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn9 net15 SE net13 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn10 net13 D net16 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn8 net16 net9 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn3 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn0 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn6 net13 ncki net3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn4 net3 cki net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.2e-07 L=6.4e-07
M_tn16_8 VSS net6 Q VPW nfet_05v0 W=8.2e-07 L=6e-07
M_tp11 net9 SE VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp10 net11 SI VDD VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp1 net8 net9 net11 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp8 net12 D net8 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp7 VDD SE net12 VNW pfet_05v0 W=6.3e-07 L=5e-07
M_tp4 ncki CLK VDD VNW pfet_05v0 W=9.25e-07 L=5e-07
M_tp0 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp9 net3 cki net8 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp6 net10 ncki net3 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp18 net5 ncki net4 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp17 net7 cki net5 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=6.25e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp14_2 VDD net6 Q VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4 D SE SETN SI CLK Q VDD VNW VPW VSS
M_tn11 net9 SE VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn7 VSS SI net15 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn9 net15 SE net13 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn10 net13 D net16 VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn8 net16 net9 VSS VPW nfet_05v0 W=3.8e-07 L=6e-07
M_tn3 ncki CLK VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn0 cki ncki VSS VPW nfet_05v0 W=4.65e-07 L=6e-07
M_tn6 net13 ncki net3 VPW nfet_05v0 W=4.75e-07 L=6e-07
M_tn4 net3 cki net14 VPW nfet_05v0 W=4.75e-07 L=6e-07
M_tn5 VSS net4 net14 VPW nfet_05v0 W=4.75e-07 L=6e-07
M_tn2 net0 net3 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn1 net4 SETN net0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn13 net5 cki net4 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn12 net7 ncki net5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_tn14 net1 SETN net7 VPW nfet_05v0 W=3.7e-07 L=6e-07
M_tn15 VSS net6 net1 VPW nfet_05v0 W=3.7e-07 L=6e-07
M_tn18 net6 net5 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn18_45 net6 net5 VSS VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_8 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_23 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tn16_8_32 VSS net6 Q VPW nfet_05v0 W=8.15e-07 L=6e-07
M_tp11 net9 SE VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp10 net11 SI VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp1 net8 net9 net11 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp8 net12 D net8 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp7 VDD SE net12 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp4 ncki CLK VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp0 cki ncki VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp9 net3 cki net8 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp6 net10 ncki net3 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp5 VDD net4 net10 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_tp3 net4 net3 VDD VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp2 VDD SETN net4 VNW pfet_05v0 W=8.15e-07 L=5e-07
M_tp18 net5 ncki net4 VNW pfet_05v0 W=4.15e-07 L=5e-07
M_tp17 net7 cki net5 VNW pfet_05v0 W=4.15e-07 L=5e-07
M_tp12 net7 SETN VDD VNW pfet_05v0 W=4.7e-07 L=5e-07
M_tp13 VDD net6 net7 VNW pfet_05v0 W=4.7e-07 L=5e-07
M_tp16 net6 net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp16_52 net6 net5 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp14_2 VDD net6 Q VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp14_18 VDD net6 Q VNW pfet_05v0 W=1.22e-06 L=5e-07
M_tp14_2_28 VDD net6 Q VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
M_n_tran_1 VSS A A VPW nfet_05v0 W=0.82U L=0.600000U
M_p_tran_2 VDD A Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
M_n_tran_1 VSS A ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_transistor_0 VDD A A VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
M_i_6 net_2 A2 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_7 VSS A1 net_2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 net_0 I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 net_0 A2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8 I A2 VDD VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_9 VDD A1 I VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_5 ZN I VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_3 net_1 A1 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_4 VDD A2 net_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
M_i_8 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_9 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_4 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VSS A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10 net_2 A2 I VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_11 VDD A1 net_2 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_7 net_1 I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5 Z_neg A1 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6 net_1 A2 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 ZN Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xnor2_4 A1 A2 ZN VDD VNW VPW VSS
M_i_8 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_9 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_4 Z_neg I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 net_0 A1 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 VSS A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 ZN Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 ZN Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS Z_neg ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10 net_2 A2 I VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_11 VDD A1 net_2 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_7 net_1 I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_5 Z_neg A1 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_6 net_1 A2 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_0 ZN Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 ZN Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_12 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_13 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 I2 I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 net_0 A1 I2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_16 net_5 I2 I3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_17 VSS A3 net_5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_8 net_2 I3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6 ZN A3 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7 net_2 I2 ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_14 net_4 A2 I VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_15 VDD A1 net_4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_5 net_1 I VDD VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_3 I2 A1 net_1 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_4 net_1 A2 I2 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_18 I3 I2 VDD VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_19 VDD A3 I3 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_11 ZN I3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_9 net_3 A3 ZN VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_10 VDD I2 net_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_14 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_15 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 I2 I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 net_0 A1 I2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_18 I3 I2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_19 VSS A3 I3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_10 Z_neg I3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8 net_2 A3 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9 VSS I2 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_1 VSS Z_neg ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_0 ZN Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_16 net_4 A2 I VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_17 VDD A1 net_4 VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_5 net_1 I VDD VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_3 I2 A1 net_1 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_4 net_1 A2 I2 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_20 net_5 I2 I3 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_21 VDD A3 net_5 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_13 net_3 I3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11 Z_neg A3 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_12 net_3 I2 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 VDD Z_neg ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 ZN Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xnor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
M_i_14 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_15 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 I2 I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 net_0 A1 I2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_18 I3 I2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_19 VSS A3 I3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_10 Z_neg I3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8 net_2 A3 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9 VSS I2 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_3 VSS Z_neg ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_2 ZN Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_1 VSS Z_neg ZN VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_0 ZN Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_16 net_4 A2 I VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_17 VDD A1 net_4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_5 net_1 I VDD VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_3 I2 A1 net_1 VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_4 net_1 A2 I2 VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_20 net_5 I2 I3 VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_21 VDD A3 net_5 VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_13 net_3 I3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_11 Z_neg A3 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_12 net_3 I2 Z_neg VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_3 VDD Z_neg ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_2 ZN Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 VDD Z_neg ZN VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 ZN Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
M_i_6 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_7 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 Z I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0 net_0 A1 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8 net_2 A2 I VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_9 VDD A1 net_2 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_5 net_1 I VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_3 Z A1 net_1 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_4 net_1 A2 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
M_i_8 net_2 A2 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_9 VSS A1 net_2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_4 net_0 I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 Z_neg A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 net_0 A2 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10 I A2 VDD VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_11 VDD A1 I VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_7 Z_neg I VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5 net_1 A1 Z_neg VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6 VDD A2 net_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
M_i_8 net_2 A2 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_9 VSS A1 net_2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_4 net_0 I VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_2 Z_neg A1 net_0 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_3 net_0 A2 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_2 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_0_3 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_10 I A2 VDD VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_11 VDD A1 I VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_7 Z_neg I VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_5 net_1 A1 Z_neg VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_6 VDD A2 net_1 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_1_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_1_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
M_i_12 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_13 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 I2 I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 net_0 A1 I2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_16 I3 I2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_17 VSS A3 I3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_8 Z I3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6 net_2 A3 Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_7 VSS I2 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_14 net_4 A2 I VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_15 VDD A1 net_4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_5 net_1 I VDD VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_3 I2 A1 net_1 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_4 net_1 A2 I2 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_18 net_5 I2 I3 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_19 VDD A3 net_5 VNW pfet_05v0 W=5.65e-07 L=5e-07
M_i_11 net_3 I3 VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_9 Z A3 net_3 VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_10 net_3 I2 Z VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
M_i_14 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_15 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 I2 I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 net_0 A1 I2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_18 net_5 I2 I3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_19 VSS A3 net_5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_10 net_2 I3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8 Z_neg A3 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9 net_2 I2 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_16 net_4 A2 I VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_17 VDD A1 net_4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_5 net_1 I VDD VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_3 I2 A1 net_1 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_4 net_1 A2 I2 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_20 I3 I2 VDD VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_21 VDD A3 I3 VNW pfet_05v0 W=5.6e-07 L=5e-07
M_i_13 Z_neg I3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11 net_3 A3 Z_neg VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_12 VDD I2 net_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__xor3_4 A1 A2 A3 Z VDD VNW VPW VSS
M_i_14 I A2 VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_15 VSS A1 I VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_2 I2 I VSS VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_0 net_0 A1 I2 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_1 VSS A2 net_0 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_18 net_5 I2 I3 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_19 VSS A3 net_5 VPW nfet_05v0 W=3.6e-07 L=6e-07
M_i_10 net_2 I3 VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_8 Z_neg A3 net_2 VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_9 net_2 I2 Z_neg VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_3 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_2 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_1 VSS Z_neg Z VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_6_0 Z Z_neg VSS VPW nfet_05v0 W=8.2e-07 L=6e-07
M_i_16 net_4 A2 I VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_17 VDD A1 net_4 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_5 net_1 I VDD VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_3 I2 A1 net_1 VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_4 net_1 A2 I2 VNW pfet_05v0 W=3.85e-07 L=5e-07
M_i_20 I3 I2 VDD VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_21 VDD A3 I3 VNW pfet_05v0 W=3.6e-07 L=5e-07
M_i_13 Z_neg I3 VDD VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_11 net_3 A3 Z_neg VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_12 VDD I2 net_3 VNW pfet_05v0 W=1.095e-06 L=5e-07
M_i_7_3 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_2 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_1 VDD Z_neg Z VNW pfet_05v0 W=1.22e-06 L=5e-07
M_i_7_0 Z Z_neg VDD VNW pfet_05v0 W=1.22e-06 L=5e-07
.ENDS


******* EOF

.END