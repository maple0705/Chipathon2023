* NGSPICE file created from user_proj_sarlogic.ext - technology: gf180mcuD

.subckt user_proj_sarlogic CLK COMP_CLK COMP_OUT DIGITAL_OUT[0] DIGITAL_OUT[1] DIGITAL_OUT[2]
+ DIGITAL_OUT[3] DIGITAL_OUT[4] DIGITAL_OUT[5] EOC XRST SC SDAC[0] SDAC[1] SDAC[2]
+ SDAC[3] SDAC[4] SDAC[5] SDAC[6] vccd1 vssd1
X0 a_25660_24328# a_25572_24372# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 vccd1 a_27116_20759# a_27028_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 SDAC[5] a_1772_20408# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_12424_13484# a_11460_13880# a_12220_13484# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 vccd1 a_22748_7080# a_22660_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 vssd1 a_8153_25200# a_8048_25244# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X6 vccd1 a_25772_17623# a_25684_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_6999_13188# a_6543_12612# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X8 a_19612_3944# a_19524_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X9 a_18853_22826# a_18733_23269# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X10 vccd1 a_5685_16533# a_6095_16532# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X11 a_15244_5079# a_15156_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 a_1692_26427# a_8153_25200# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X13 a_4264_17020# a_2052_17016# a_3324_16576# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X14 a_24640_25940# a_24004_22804# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X15 a_6527_24047# a_5627_23544# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
D0 vssd1 a_1804_21723# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X16 a_18268_11784# a_18180_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X17 vssd1 a_5084_25560# a_13216_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X18 vssd1 a_20196_25940# a_21392_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X19 vccd1 a_19544_24416# a_19352_24460# vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X20 vccd1 a_27116_14487# a_27028_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X21 a_10316_6647# a_10228_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X22 a_2016_19739# a_1604_20152# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_25660_18056# a_25572_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X24 a_1692_18528# a_6440_18056# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X25 a_19477_18100# a_19357_18632# a_18733_18565# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X26 a_1892_14180# a_1772_14136# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X27 vccd1 a_27116_11351# a_27028_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X28 a_25660_14920# a_25572_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X29 vssd1 a_6266_14756# a_6742_14180# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X30 vccd1 a_2588_5512# a_2500_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X31 a_8583_20856# a_8736_25940# a_7452_21280# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X32 vccd1 a_23084_9783# a_22996_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X33 a_6118_10836# a_5642_10260# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X34 a_1892_11044# a_1772_11000# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X35 a_22448_22424# a_21684_22020# a_22244_22424# vccd1 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X36 a_3816_15452# a_2016_15035# a_2876_15008# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X37 vccd1 a_8300_5079# a_8212_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X38 a_28012_6647# a_27924_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X39 vccd1 a_15692_8215# a_15604_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D1 a_2444_24328# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X40 vssd1 a_1772_12568# SDAC[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X41 vccd1 a_23084_6647# a_22996_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X42 a_12560_16976# a_11548_13824# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X43 a_16588_14487# a_16500_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X44 vccd1 a_13672_13884# a_14089_13744# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X45 a_10192_8692# a_7988_3608# vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X46 vccd1 a_10452_18840# a_8736_19363# vccd1 pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X47 a_24540_16488# a_24452_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X48 vccd1 a_17585_20856# a_9263_20408# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X49 a_1692_10688# a_6328_17342# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X50 DIGITAL_OUT[2] a_17024_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X51 a_7190_18884# a_6358_19378# a_7042_19460# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X52 vccd1 a_24204_18056# a_24116_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X53 a_19948_17623# a_19860_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X54 vccd1 a_4041_24812# a_3981_24460# vccd1 pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X55 vccd1 a_16520_20128# a_6388_6390# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X56 a_8968_11132# a_8040_11503# a_8800_11132# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X57 vssd1 a_11961_12656# a_11856_12700# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X58 a_12668_5512# a_12580_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X59 a_22748_19624# a_22660_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X60 vssd1 a_7302_10836# a_7778_10835# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X61 a_14860_20807# a_14552_20856# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X62 a_24316_21192# a_24228_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X63 vccd1 a_25660_8648# a_25572_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D2 a_2140_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X64 vccd1 a_26332_3511# a_26244_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X65 DIGITAL_OUT[1] a_13216_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X66 vccd1 a_25660_5512# a_25572_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X67 a_4348_7909# a_5577_9040# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X68 vccd1 a_26556_10216# a_26468_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X69 a_18604_11351# a_18516_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X70 a_5084_25560# a_4628_25248# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X71 a_6571_17108# a_6095_16532# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X72 a_17820_8648# a_17732_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X73 a_7302_10836# a_6470_10260# a_7154_10260# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X74 a_7706_22424# a_5836_22760# a_1916_22021# vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X75 a_13452_9783# a_13364_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X76 a_5836_22760# a_14649_21584# vssd1 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X77 vccd1 a_18716_16488# a_18628_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X78 a_14068_23992# a_13508_23588# a_13940_23588# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X79 a_3036_8215# a_2948_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X80 SDAC[2] a_1772_9432# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X81 vccd1 a_27564_23895# a_27476_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X82 vssd1 a_14392_14181# a_8335_13352# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X83 vccd1 a_14460_7080# a_14372_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X84 vssd1 a_12579_24765# a_8492_24328# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X85 a_11544_12700# a_9332_12695# a_10604_12967# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X86 vccd1 a_27564_20759# a_27476_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X87 a_22636_20759# a_22548_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X88 a_11548_3511# a_11460_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X89 vccd1 a_8519_13836# a_8721_14920# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X90 vccd1 a_1772_9432# SDAC[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X91 a_11799_16488# a_12560_16976# a_12351_16620# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X92 DIGITAL_OUT[3] a_18256_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X93 a_10901_24142# a_10781_23544# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X94 a_22188_12919# a_22100_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X95 vccd1 a_1772_6296# SDAC[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X96 vccd1 a_13533_24904# a_13653_24372# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X97 DIGITAL_OUT[0] a_9408_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X98 EOC a_25648_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X99 a_19724_5079# a_19636_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X100 vccd1 a_1772_3160# SDAC[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X101 a_5276_5512# a_5188_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X102 vccd1 a_17859_24373# a_19760_23992# vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X103 vssd1 a_5836_22760# a_4631_20408# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X104 vssd1 a_3564_25112# a_1772_25112# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X105 vssd1 a_20196_25940# a_21392_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X106 a_21852_3944# a_21764_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X107 a_5936_25560# a_5524_25239# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X108 vccd1 a_27564_14487# a_27476_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X109 a_22636_14487# a_22548_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X110 a_9408_25940# a_2052_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X111 a_1692_18528# a_6440_18056# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X112 a_22636_11351# a_22548_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X113 vccd1 a_27564_11351# a_27476_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X114 a_11405_23544# a_2672_21782# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X115 vccd1 a_27564_9783# a_27476_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X116 vccd1 a_16364_11351# a_16276_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X117 vccd1 a_1772_23544# SDAC[6] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X118 vccd1 a_27564_6647# a_27476_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X119 vccd1 a_1772_20408# SDAC[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X120 a_1772_20408# a_3564_20408# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X121 vccd1 a_22748_16488# a_22660_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X122 a_2140_7080# a_2052_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X123 a_9076_15704# a_5019_20408# a_13780_18884# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X124 a_3619_17272# a_3949_17272# a_4069_17870# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X125 a_8524_5512# a_8436_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X126 vccd1 a_14348_5079# a_14260_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X127 vccd1 a_28012_17623# a_27924_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X128 a_3619_14136# a_3949_14136# a_4069_14734# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X129 vccd1 a_22636_8215# a_22548_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X130 a_10372_24372# a_9900_24756# a_10224_24372# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X131 a_19357_23336# a_10732_24328# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
D3 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X132 vccd1 a_6383_21028# a_6839_21006# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X133 a_12880_13884# a_12732_13440# a_12712_13884# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X134 vccd1 a_20396_20759# a_20308_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X135 a_2772_19756# a_1604_20152# a_2568_19756# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X136 a_8156_17584# a_9800_18056# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X137 a_8636_7080# a_8548_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X138 a_4481_24757# a_10192_8692# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X139 vccd1 a_21404_10216# a_21316_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X140 a_13126_12404# a_12650_11828# a_12854_11828# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X141 a_8132_24372# a_2444_24328# a_7984_24372# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X142 vccd1 a_9900_24756# a_9812_24856# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X143 a_4752_15704# a_5020_15796# vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X144 COMP_CLK a_2444_26249# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X145 a_26220_23895# a_26132_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X146 a_2116_14584# a_1996_11000# a_1872_14602# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X147 a_7605_13396# a_7485_13928# a_6861_13861# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X148 a_10111_17775# a_9211_17272# vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X149 a_18268_3944# a_18180_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X150 a_2116_11448# a_1996_11000# a_1872_11466# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X151 vccd1 a_13564_3944# a_13476_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X152 a_15244_8648# a_15156_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X153 a_12502_12404# a_12026_11828# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X154 a_13999_22596# a_13375_22020# a_13831_22596# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X155 a_7167_13188# a_6543_12612# a_6999_13188# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X156 vccd1 a_22412_23895# a_22324_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D4 a_5940_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X157 a_2856_23292# a_2016_22875# a_2568_22892# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
D5 vssd1 a_2220_24686# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X158 a_17932_9783# a_17844_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X159 a_25100_25463# a_25012_25560# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X160 a_17632_21976# a_16388_22424# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X161 a_5836_22760# a_14649_21584# vssd1 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X162 a_2856_20156# a_2016_19739# a_2568_19756# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X163 vssd1 a_15848_20128# a_3564_20408# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X164 vccd1 a_20396_11351# a_20308_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X165 a_14840_20540# a_14000_20856# a_14552_20856# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X166 vccd1 a_6531_13789# a_6239_12568# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X167 a_27317_24372# a_27197_24904# a_26573_24837# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X168 vssd1 a_1772_9432# SDAC[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X169 a_2364_15052# a_2264_15008# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X170 a_14089_13744# a_13672_13884# a_14465_13884# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X171 a_2364_19756# a_1792_16532# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X172 a_27900_13352# a_27812_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X173 a_6266_10260# a_5642_10260# a_6118_10836# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X174 vssd1 a_8736_19363# a_9476_17016# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X175 vccd1 a_9980_3944# a_9892_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X176 vccd1 a_21404_7080# a_21316_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X177 vccd1 a_17820_10216# a_17732_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X178 a_27900_10216# a_27812_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X179 vssd1 a_13686_12404# a_14162_12403# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X180 EOC a_25648_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X181 vccd1 a_4481_24757# a_4041_24812# vccd1 pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X182 vccd1 a_26243_24765# a_22604_21976# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X183 vccd1 a_4403_21582# a_4315_21237# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.6561p ps=3.51u w=1.215u l=0.5u
X184 vssd1 a_4236_26254# a_2444_26249# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X185 a_12375_14964# a_11919_14964# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X186 vccd1 a_23868_22327# a_23780_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X187 vccd1 a_6172_3944# a_6084_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X188 a_19164_19191# a_19076_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X189 a_1772_9432# a_3564_9432# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X190 a_8232_11390# a_7639_11459# a_8968_11132# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X191 a_9408_25940# a_2052_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X192 vccd1 a_12332_5079# a_12244_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X193 a_1772_6296# a_3564_6296# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X194 vccd1 a_20620_8215# a_20532_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X195 a_3999_21676# a_4233_23152# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X196 vccd1 a_1772_23544# SDAC[6] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X197 a_12337_12700# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X198 a_15692_5079# a_15604_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X199 a_1772_3160# a_3564_3160# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X200 a_22748_8648# a_22660_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X201 DIGITAL_OUT[4] a_21392_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X202 a_12581_14136# a_8435_13397# a_13364_12612# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X203 vccd1 a_1772_20408# SDAC[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D6 vssd1 a_2140_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X204 a_2444_24328# a_5836_22760# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
D7 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X205 a_1692_17302# a_10900_14964# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X206 a_10903_10216# a_11559_10304# a_11455_10348# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X207 a_21616_25560# a_21204_25239# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X208 a_7988_19668# a_7540_20199# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X209 a_6328_17342# a_8156_17584# vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X210 vccd1 a_18828_5079# a_18740_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X211 a_10764_6647# a_10676_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X212 a_12533_9476# a_12413_9432# a_11789_9432# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X213 a_4573_11000# a_1872_11466# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X214 a_16388_25940# a_15940_26471# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X215 a_17221_20453# a_16217_20496# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X216 a_16252_3944# a_16164_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X217 vssd1 a_11628_18056# a_13776_18100# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X218 a_14188_18884# a_5019_20408# a_9076_15704# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X219 vssd1 a_1804_21723# a_4516_9521# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X220 a_4569_12176# a_4152_12316# a_4945_12316# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X221 vccd1 a_21852_10216# a_21764_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X222 vccd1 a_26108_14920# a_26020_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X223 vccd1 a_1692_18528# a_1604_20152# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X224 a_11324_5512# a_11236_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X225 a_6971_9176# a_3479_18840# a_1772_14136# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X226 vccd1 a_26108_11784# a_26020_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X227 vccd1 a_4681_16880# a_4576_17020# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X228 a_12628_13484# a_11460_13880# a_12424_13484# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X229 vccd1 a_17024_25940# DIGITAL_OUT[2] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X230 a_22771_24765# a_23101_24837# a_23221_24947# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X231 vccd1 a_5836_22760# a_9956_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X232 a_14649_21584# a_14232_21724# a_15025_21724# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X233 a_14860_20807# a_14552_20856# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
D8 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X234 vccd1 a_22860_23895# a_22772_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X235 a_5972_17720# a_5524_17361# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X236 vccd1 a_17036_8215# a_16948_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D9 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X237 a_19276_14487# a_19188_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X238 vccd1 a_20508_3944# a_20420_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X239 vssd1 a_15849_22804# a_16192_25244# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X240 vssd1 CLK a_13496_17337# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X241 vccd1 a_4481_24757# a_11787_20027# vccd1 pfet_06v0 ad=0.33755p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X242 a_4128_15452# a_2016_15035# a_3816_15452# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X243 a_6235_26516# a_5759_25940# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X244 vccd1 a_26780_3511# a_26692_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X245 a_10204_3511# a_10116_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X246 a_13686_12404# a_12854_11828# a_13538_11828# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X247 a_7932_20453# a_3703_18840# a_8433_20152# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X248 a_9659_9176# a_8121_13016# a_7852_9006# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X249 a_27004_21192# a_26916_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X250 vccd1 a_21292_17623# a_21204_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X251 a_10452_18840# a_16744_22042# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X252 vccd1 a_7224_23934# a_7032_24047# vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X253 vccd1 a_14232_21724# a_14649_21584# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
D10 vssd1 a_1804_21723# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X254 vccd1 a_27004_8648# a_26916_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X255 vssd1 a_15064_25502# a_14872_25615# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X256 vccd1 a_11628_18056# a_13776_18100# vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X257 vccd1 a_19612_7080# a_19524_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X258 a_1772_9432# a_3564_9432# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X259 SDAC[4] a_1772_15704# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X260 vccd1 a_27004_5512# a_26916_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X261 a_9868_6647# a_9780_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X262 a_11996_3511# a_11908_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X263 vccd1 a_24428_19191# a_24340_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X264 a_18716_14920# a_18628_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X265 a_28012_8215# a_27924_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X266 vssd1 a_8009_11828# a_9360_11132# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X267 vccd1 a_21740_16055# a_21652_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X268 vssd1 a_1692_17302# a_14092_14920# vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X269 a_2968_17317# a_3228_17317# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X270 vccd1 a_21740_12919# a_21652_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X271 a_4074_22020# a_3954_21976# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X272 vssd1 a_9532_19624# a_10866_20152# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X273 vccd1 a_5724_5512# a_5636_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X274 vssd1 a_16744_22042# a_10452_18840# vssd1 nfet_06v0 ad=0.151p pd=1.185u as=0.1261p ps=1.005u w=0.485u l=0.6u
X275 a_25324_20759# a_25236_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X276 vccd1 a_26220_9783# a_26132_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X277 a_13608_19712# a_13015_19712# a_14344_20156# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X278 a_2016_18171# a_1604_18584# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X279 vccd1 a_8009_11828# a_9360_11132# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X280 a_27004_11784# a_26916_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X281 a_2016_15035# a_1604_15448# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X282 vccd1 a_26220_6647# a_26132_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X283 a_9920_20096# a_11787_20027# vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X284 a_11628_18056# a_13496_17337# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X285 vssd1 a_10396_16488# a_10348_17016# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X286 vccd1 a_13776_18100# a_14708_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X287 a_20060_16488# a_19972_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X288 a_1772_14136# a_3479_18840# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X289 a_16588_9783# a_16500_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X290 DIGITAL_OUT[5] a_24640_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X291 vccd1 a_23868_21192# a_23780_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X292 a_26668_17623# a_26580_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X293 a_22636_5079# a_22548_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X294 a_12668_7080# a_12580_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X295 vccd1 a_13216_25940# DIGITAL_OUT[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X296 SC a_1772_25112# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X297 a_18604_16055# a_18516_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X298 a_19056_24816# a_12108_21664# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X299 vccd1 a_26108_22327# a_26020_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X300 a_11799_16488# a_12455_16576# a_12351_16620# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X301 vccd1 a_26556_14920# a_26468_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X302 vccd1 a_1916_17302# a_8736_19363# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X303 a_1812_17353# a_2140_17302# vssd1 vssd1 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X304 a_25324_14487# a_25236_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X305 a_15804_5512# a_15716_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X306 vccd1 a_26556_11784# a_26468_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X307 a_2876_18144# a_2568_18188# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X308 a_4464_12316# a_1940_12312# a_4152_12316# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X309 a_7175_24856# a_4815_20408# a_6991_24856# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X310 a_13776_18100# a_11628_18056# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X311 vccd1 a_14796_5079# a_14708_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X312 a_25324_11351# a_25236_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X313 vccd1 a_15356_11784# a_15268_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X314 vssd1 a_9408_25940# DIGITAL_OUT[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X315 a_21336_23589# a_5539_23589# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X316 a_9308_3511# a_9220_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D11 a_1692_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X317 a_14124_11351# a_14036_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X318 vccd1 a_19052_11351# a_18964_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X319 vccd1 a_12220_3944# a_12132_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X320 a_22748_14920# a_22660_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X321 a_4481_24757# a_10192_8692# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X322 a_10612_22892# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X323 a_7852_9006# a_8121_13016# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X324 a_8940_21590# a_4631_20408# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X325 SDAC[4] a_1772_15704# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X326 vccd1 a_3816_10748# a_4233_10608# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X327 SDAC[3] a_1772_12568# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X328 a_2052_25940# a_1604_26471# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X329 a_12073_23152# a_11656_23292# a_12449_23292# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X330 a_17585_20856# a_2220_24686# a_17605_20452# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X331 a_5600_18101# a_4672_12657# a_5412_18101# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X332 vccd1 a_18716_3944# a_18628_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X333 a_6991_24856# a_5836_22760# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X334 vccd1 a_23084_20759# a_22996_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X335 a_15692_8648# a_15604_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X336 a_21392_25940# a_20196_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X337 a_10451_23544# a_10781_23544# a_10901_24142# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X338 a_11548_13824# a_13496_15774# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X339 a_27452_21192# a_27364_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X340 vccd1 a_5836_22760# a_8736_19363# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X341 a_5817_24800# a_4913_24860# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X342 a_2672_21237# a_1916_22021# vccd1 vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X343 a_22636_19191# a_22548_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X344 vccd1 a_3619_14136# a_2264_13440# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X345 a_9920_11828# a_6388_6390# vccd1 vccd1 pfet_06v0 ad=0.224p pd=1.36u as=0.389p ps=2.02u w=0.56u l=0.5u
X346 a_22636_16055# a_22548_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X347 vccd1 a_3619_11000# a_2264_10304# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X348 a_16324_23992# a_15156_23671# a_16120_23992# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X349 a_9444_19668# a_7259_24800# a_10040_20152# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X350 a_10808_13396# a_10136_13396# vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X351 a_17372_13352# a_17284_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X352 vssd1 a_1772_23544# SDAC[6] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X353 vccd1 a_23084_14487# a_22996_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X354 a_11076_24372# a_10372_24372# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X355 vccd1 a_24876_19191# a_24788_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X356 a_7829_7908# a_7709_7864# a_7085_7864# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X357 a_17372_10216# a_17284_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X358 a_8454_21572# a_8940_21590# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X359 vccd1 a_23084_11351# a_22996_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X360 a_27900_19624# a_27812_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X361 vccd1 a_11544_12700# a_11961_12656# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X362 vccd1 a_21852_7080# a_21764_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D12 vssd1 a_1692_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X363 a_6887_22804# a_6431_22804# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X364 a_12100_22020# a_9076_15704# a_12308_22020# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X365 a_20620_5079# a_20532_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X366 a_25772_20759# a_25684_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X367 a_12359_19624# a_13015_19712# a_12911_19756# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X368 vssd1 a_3564_9432# a_1772_9432# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X369 a_8836_24372# a_8132_24372# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X370 a_21404_8648# a_21316_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X371 a_27452_11784# a_27364_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X372 a_20196_25940# a_19748_26471# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X373 a_3404_24812# a_5612_23118# a_5524_23288# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X374 a_15371_23379# a_14895_22804# a_15119_22826# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X375 vccd1 a_21404_14920# a_21316_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X376 a_11685_14734# a_11565_14136# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X377 a_16252_11784# a_16164_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X378 vccd1 a_4481_24757# a_17947_24328# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X379 vssd1 a_7259_24800# a_7628_20155# vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X380 a_11628_18056# a_13496_17337# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X381 DIGITAL_OUT[5] a_24640_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X382 vccd1 a_18984_22021# a_3564_23544# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X383 vccd1 a_21404_11784# a_21316_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X384 a_17499_24856# a_5612_23118# a_10104_22848# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X385 vccd1 a_12780_5079# a_12692_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X386 vccd1 a_13216_25940# DIGITAL_OUT[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X387 a_20620_18056# a_20532_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X388 vccd1 a_20172_18056# a_20084_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X389 a_9559_17540# a_10215_17731# a_10111_17775# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X390 vccd1 a_1692_8648# a_1604_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X391 vccd1 a_17844_25560# a_18256_25560# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X392 a_1772_15704# a_3564_15704# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X393 vccd1 a_1692_5512# a_1604_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X394 vssd1 a_1692_10688# a_6532_9559# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X395 vccd1 a_1692_17302# a_9532_19624# vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X396 vccd1 a_26556_22327# a_26468_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X397 a_25772_14487# a_25684_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X398 vssd1 a_7224_23934# a_7032_24047# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X399 a_6440_18056# a_8156_17584# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X400 a_19357_18632# a_5020_15796# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X401 a_25772_11351# a_25684_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X402 vssd1 a_9408_25940# DIGITAL_OUT[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X403 vccd1 a_9920_20096# a_13375_22020# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X404 a_14572_11351# a_14484_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X405 vccd1 a_16700_3944# a_16612_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X406 vccd1 a_18268_7080# a_18180_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X407 vccd1 a_27900_22760# a_27812_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X408 a_17036_5079# a_16948_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X409 a_6736_23632# a_1692_18528# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X410 a_8040_11503# a_7639_11459# a_6983_11268# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X411 a_28012_24328# a_27924_24372# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X412 a_15008_20540# a_14860_20807# a_14840_20540# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X413 COMP_CLK a_2444_26249# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X414 a_8736_25940# a_2500_22020# vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X415 a_14428_23544# a_17785_23632# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X416 a_11772_5512# a_11684_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X417 vccd1 a_26108_21192# a_26020_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X418 vccd1 a_4815_20408# a_4731_20872# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X419 vccd1 a_17820_14920# a_17732_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X420 vccd1 a_18380_12919# a_18292_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X421 a_12108_6647# a_12020_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X422 a_1772_25112# a_3564_25112# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X423 a_15816_23822# a_15119_24394# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X424 vccd1 a_11656_23292# a_12073_23152# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X425 vccd1 a_17820_11784# a_17732_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X426 a_11968_23292# a_9444_23288# a_11656_23292# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X427 a_2856_18588# a_2016_18171# a_2568_18188# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X428 vccd1 a_24540_10216# a_24452_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X429 a_3542_22242# a_3954_21976# a_4074_22020# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X430 vccd1 a_9900_13396# a_9532_19624# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X431 vccd1 a_17484_8215# a_17396_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X432 vccd1 a_8744_9564# a_9161_9520# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X433 vssd1 a_11664_10704# a_11559_10304# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X434 a_3703_18840# a_8454_21572# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X435 vccd1 a_27900_16488# a_27812_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X436 DIGITAL_OUT[3] a_18256_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X437 vccd1 a_20956_3944# a_20868_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X438 a_14895_24372# a_14271_24372# a_14727_24372# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X439 a_9771_22020# a_9295_22596# a_9519_22020# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X440 a_12132_19288# a_5237_19669# a_2892_18840# vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X441 vssd1 a_5076_23992# a_2892_18840# vssd1 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X442 a_4573_14136# a_4965_14136# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X443 a_2140_8215# a_2052_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X444 SDAC[2] a_1772_9432# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X445 vccd1 a_8940_21590# a_10599_11829# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X446 vssd1 a_1772_23544# SDAC[6] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X447 vccd1 a_8736_19363# a_9476_17016# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X448 a_8524_6647# a_8436_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X449 a_6563_11784# a_1996_11000# a_7524_8692# vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X450 a_6747_22020# a_6271_22596# a_6495_22020# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X451 a_4573_11000# a_1872_11466# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X452 a_22300_11784# a_22212_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X453 a_15456_19368# a_14708_18100# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X454 a_1772_15704# a_3564_15704# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X455 a_10652_3511# a_10564_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X456 vccd1 a_7628_5512# a_7540_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X457 DIGITAL_OUT[2] a_17024_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X458 a_3728_24460# a_2724_24856# a_3524_24460# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X459 a_19477_21812# a_19357_21768# a_18733_21701# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X460 a_14796_10216# a_14708_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X461 a_12100_22020# a_12860_21976# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X462 a_1692_18528# a_6440_18056# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X463 a_1772_12568# a_3564_12568# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X464 a_20172_12919# a_20084_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X465 vccd1 a_27452_8648# a_27364_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X466 a_11872_13467# a_11460_13880# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X467 vccd1 a_4236_26254# a_2444_26249# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X468 a_26693_24394# a_26573_24837# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X469 a_18853_21811# a_18733_21701# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X470 vccd1 a_19948_16055# a_19860_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X471 a_13494_14136# a_8519_13836# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X472 vccd1 a_27452_5512# a_27364_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X473 a_4380_5512# a_4292_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X474 SC a_1772_25112# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X475 vccd1 a_15849_22804# a_16192_25244# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X476 vssd1 a_7485_15496# a_7605_15540# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X477 vccd1 a_1692_18885# a_4628_23633# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X478 a_23845_24948# a_23725_24904# a_23101_24837# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X479 vccd1 a_1804_21723# a_1716_21767# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X480 a_5895_21372# a_5547_21551# a_4771_21192# vssd1 nfet_06v0 ad=0.1989p pd=1.465u as=93.59999f ps=0.88u w=0.36u l=0.6u
X481 vccd1 a_9800_18056# a_8156_17584# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X482 vccd1 a_21852_14920# a_21764_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X483 a_20620_14487# a_20532_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X484 a_4609_13884# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X485 a_19612_8648# a_19524_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X486 a_6944_9880# a_6532_9559# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X487 vccd1 a_21852_11784# a_21764_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X488 a_13900_6647# a_13812_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X489 EOC a_25648_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X490 a_11324_7080# a_11236_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X491 a_15244_9783# a_15156_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X492 a_4609_10748# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X493 a_12732_13440# a_12424_13484# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X494 vccd1 a_6844_3511# a_6756_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X495 a_18268_16488# a_18180_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X496 vccd1 a_16252_7080# a_16164_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X497 a_6440_18056# a_8156_17584# vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X498 vccd1 a_16217_20496# a_16112_20540# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X499 vccd1 a_27116_19191# a_27028_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X500 vccd1 a_10320_17360# a_10215_17731# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X501 vccd1 a_7001_19668# a_2264_22848# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X502 a_2544_19306# a_2444_18840# vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X503 a_16428_23943# a_16120_23992# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X504 vccd1 a_13452_5079# a_13364_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X505 a_28012_20759# a_27924_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X506 a_4128_20156# a_2016_19739# a_3816_20156# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X507 a_6907_12404# a_6431_11828# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X508 vccd1 a_21740_8215# a_21652_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X509 vccd1 a_19556_23992# a_20260_23588# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X510 a_18256_25560# a_17844_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X511 a_14176_20156# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X512 vccd1 a_14428_23544# a_17396_25201# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X513 vccd1 a_4481_24757# a_19804_24460# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X514 vccd1 a_26556_21192# a_26468_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X515 a_23644_3944# a_23556_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X516 a_2116_24856# a_1996_24328# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X517 vssd1 a_18403_23197# a_13820_23544# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X518 a_9756_3511# a_9668_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X519 a_7988_3608# a_7540_3249# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X520 a_17372_3944# a_17284_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X521 vccd1 a_10192_8692# a_4481_24757# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X522 a_28012_14487# a_27924_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X523 a_1804_21723# a_12132_26424# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X524 a_13686_12404# a_12854_11828# a_13518_12404# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X525 a_4128_15452# a_1604_15448# a_3816_15452# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X526 a_28012_11351# a_27924_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X527 vccd1 a_15916_11351# a_15828_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X528 a_7301_7608# a_1692_17302# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X529 a_13216_25940# a_5084_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X530 vssd1 a_6328_17342# a_1692_10688# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X531 a_1916_17302# a_13494_14136# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X532 vccd1 a_24428_8215# a_24340_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X533 a_17585_20856# a_2052_19288# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X534 a_2876_15008# a_2568_15052# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X535 a_10500_25560# a_9332_25239# a_10296_25560# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X536 a_8617_15448# a_4492_18840# a_8433_15448# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X537 a_8624_14602# a_8519_13836# a_8644_14181# vssd1 nfet_06v0 ad=0.4137p pd=1.9u as=0.2119p ps=1.335u w=0.815u l=0.6u
X538 vccd1 a_11760_11828# a_13280_10748# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X539 vccd1 a_1916_17302# a_8852_15704# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X540 a_7960_23676# a_7032_24047# a_7792_23676# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X541 vccd1 a_6060_5079# a_5972_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X542 vccd1 a_14908_3511# a_14820_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X543 a_14895_22804# a_14271_22804# a_14747_23380# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X544 a_15351_22826# a_14895_22804# a_15119_22826# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X545 SDAC[3] a_1772_12568# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X546 vccd1 a_12413_9432# a_12533_10052# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X547 vccd1 a_15356_3944# a_15268_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X548 vccd1 a_27004_18056# a_26916_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X549 a_10036_16532# a_9476_17016# a_9908_17016# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X550 vssd1 a_1692_17302# a_10532_15448# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1148p ps=1.1u w=0.82u l=0.6u
X551 a_1916_17302# a_13494_14136# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X552 a_7672_20453# a_7932_20453# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X553 a_5860_14964# a_5412_15495# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X554 vccd1 a_9800_18056# a_8156_17584# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X555 a_10408_22892# a_9444_23288# a_10204_22892# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X556 vssd1 a_4481_24757# a_15008_20540# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X557 a_25324_19191# a_25236_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X558 a_22188_17623# a_22100_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X559 vssd1 a_9900_24756# a_13508_23588# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X560 a_7717_15748# a_7597_15704# a_6973_15704# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X561 vccd1 a_10428_5512# a_10340_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X562 vssd1 a_4681_16880# a_4576_17020# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X563 a_25324_16055# a_25236_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X564 a_15804_7080# a_15716_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X565 a_19724_9783# a_19636_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X566 a_10612_22892# a_9444_23288# a_10408_22892# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X567 a_10500_13016# a_9332_12695# a_10296_13016# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X568 a_2672_21237# a_3004_21664# a_2672_21782# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X569 vccd1 a_27564_19191# a_27476_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X570 a_21852_8648# a_21764_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X571 vccd1 a_4815_20408# a_8736_19363# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X572 vssd1 a_7167_13188# a_7643_12612# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X573 vccd1 a_12579_24765# a_8492_24328# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X574 vssd1 a_5685_16533# a_6095_16532# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X575 vccd1 a_3816_15452# a_4233_15312# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X576 vccd1 a_17932_5079# a_17844_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X577 vccd1 a_12108_21664# a_15156_23671# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X578 vccd1 a_8764_15749# a_10228_15793# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X579 a_8752_8648# a_9161_9520# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X580 a_1772_25112# a_3564_25112# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X581 a_7225_22424# a_6495_22020# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X582 a_3912_8780# a_3360_8763# a_3708_8780# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X583 a_4716_25204# a_11961_25200# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X584 vssd1 a_1772_20408# SDAC[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X585 a_17024_25940# a_16388_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X586 a_10575_21720# a_2220_24686# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X587 a_9076_15704# a_4815_20408# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X588 a_11961_25200# a_11544_25244# a_12337_25244# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X589 vssd1 a_23833_25200# a_23728_25244# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X590 a_10204_22892# a_10104_22848# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X591 a_6271_22596# a_5647_22020# a_6123_22020# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X592 vccd1 a_10452_18840# a_8736_19363# vccd1 pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X593 a_18716_19191# a_18628_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X594 a_3024_13884# a_2876_13440# a_2856_13884# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X595 vccd1 a_3036_5512# a_2948_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X596 a_24316_22327# a_24228_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X597 a_17484_5079# a_17396_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X598 a_10244_24856# a_8492_24328# vssd1 vssd1 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X599 a_22277_22804# a_22157_23336# a_21533_23269# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X600 a_10584_22042# a_9444_19668# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.151p ps=1.185u w=0.36u l=0.6u
X601 vccd1 CLK a_13496_17337# vccd1 pfet_06v0 ad=0.3608p pd=2.52u as=0.2542p ps=1.44u w=0.82u l=0.5u
X602 a_11628_18056# a_13496_17337# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X603 vccd1 a_16140_8215# a_16052_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X604 a_3024_10748# a_2876_10304# a_2856_10748# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X605 vssd1 a_24004_22804# a_24640_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X606 vccd1 a_5817_24800# a_5137_24860# vccd1 pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X607 a_6692_25560# a_5524_25239# a_6488_25560# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X608 a_23644_23291# a_23833_25200# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X609 a_15916_23992# a_15816_23822# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X610 a_18268_8648# a_18180_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X611 a_13216_25940# a_5084_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X612 a_4180_18884# a_4672_12657# a_2220_14136# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X613 a_24092_13352# a_24004_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X614 a_12556_6647# a_12468_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X615 a_17260_11351# a_17172_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X616 a_21203_23197# a_21533_23269# a_21653_23379# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X617 a_3479_18840# a_6943_16554# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X618 a_1872_14602# a_1996_11000# a_1892_14180# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X619 a_24092_10216# a_24004_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X620 a_16324_23992# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X621 a_26108_22760# a_26020_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X622 a_1872_11466# a_1996_11000# a_1892_11044# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X623 vccd1 a_17372_16488# a_17284_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X624 a_1772_12568# a_3564_12568# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X625 a_5795_21280# a_1692_18528# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X626 vssd1 a_13496_17337# a_11628_18056# vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X627 a_13116_5512# a_13028_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X628 a_15849_22804# a_15119_22826# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X629 a_21292_20759# a_21204_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X630 a_6531_13789# a_6861_13861# a_6981_13418# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X631 a_7224_23934# a_6736_23632# a_7484_23992# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X632 a_12499_20152# a_12359_19624# a_11787_20027# vssd1 nfet_06v0 ad=0.217p pd=1.515u as=0.3586p ps=2.51u w=0.815u l=0.6u
X633 vssd1 a_11548_13824# a_13588_20535# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X634 a_27900_18056# a_27812_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X635 vccd1 a_27452_18056# a_27364_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X636 vccd1 a_13497_14964# a_14176_17020# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X637 vssd1 a_5544_7584# a_3564_12568# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X638 a_8048_25244# a_5936_25560# a_7736_25244# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X639 vccd1 a_5836_22760# a_8736_19363# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X640 a_8972_6647# a_8884_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X641 a_27900_14920# a_27812_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X642 a_5137_24860# a_2724_24856# a_4913_24860# vssd1 nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X643 a_14403_24328# a_14068_23992# vccd1 vccd1 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X644 a_15804_3511# a_15716_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X645 a_25772_19191# a_25684_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X646 a_5600_18101# a_1692_17302# a_5620_18584# vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X647 vccd1 a_14908_5512# a_14820_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X648 a_6284_25560# a_2096_24372# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X649 a_8529_25244# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X650 a_25772_16055# a_25684_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X651 a_18403_23197# a_18733_23269# a_18853_22826# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X652 vssd1 a_2444_26249# COMP_CLK vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X653 a_10451_23544# a_10781_23544# a_10901_23588# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
D13 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X654 a_18828_14487# a_18740_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X655 vccd1 a_5500_3511# a_5412_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X656 a_9532_5512# a_9444_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X657 a_21292_14487# a_21204_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X658 vssd1 a_12158_11784# a_12026_11828# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X659 a_5936_25560# a_5524_25239# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X660 a_15064_25502# a_14471_25571# a_15800_25244# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X661 a_12309_14756# a_12189_14136# a_11565_14136# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X662 a_4116_8780# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X663 a_21292_11351# a_21204_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X664 a_16388_22424# a_15940_22065# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X665 vccd1 a_19357_18632# a_19477_18100# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X666 a_4609_23292# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X667 a_11032_13880# a_8721_14920# a_10808_13880# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X668 a_15692_9783# a_15604_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X669 vssd1 a_14649_21584# a_5836_22760# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X670 a_16593_20540# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X671 a_4609_20156# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X672 a_11936_17404# a_10215_17731# a_10808_17662# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X673 vccd1 a_9612_15704# a_8764_15749# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4012p ps=1.85u w=1.13u l=0.5u
X674 a_21740_5079# a_21652_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X675 a_11772_7080# a_11684_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X676 vccd1 a_24092_8648# a_24004_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X677 a_14708_18100# a_13776_18100# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X678 vccd1 a_24540_14920# a_24452_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X679 a_8863_13880# a_8437_10291# a_8435_13397# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X680 vccd1 a_24092_5512# a_24004_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X681 a_7348_21324# a_5547_21551# a_6499_21264# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.19315p ps=1.27u w=0.505u l=0.5u
X682 a_4088_7909# a_4348_7909# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X683 vccd1 a_24540_11784# a_24452_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X684 a_22300_3944# a_22212_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X685 vssd1 a_18256_25560# DIGITAL_OUT[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X686 a_4233_13744# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X687 vccd1 a_10316_6647# a_10228_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X688 vccd1 a_20060_10216# a_19972_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X689 a_13533_24904# a_4716_25204# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X690 vccd1 a_26108_19624# a_26020_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X691 vccd1 a_25648_25560# EOC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X692 a_24764_22327# a_24676_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X693 vccd1 a_28012_9783# a_27924_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X694 a_9920_20096# a_11787_20027# vssd1 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X695 vccd1 a_28012_6647# a_27924_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D14 a_6388_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X696 a_5831_11000# a_7526_10282# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X697 vccd1 a_14403_24328# a_14271_24372# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X698 vccd1 a_4684_7564# a_2600_11872# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X699 a_24428_5079# a_24340_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X700 vccd1 a_16588_14487# a_16500_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X701 a_15064_12613# a_14350_13016# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X702 a_6702_10260# a_6266_10260# a_6470_10260# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X703 a_11068_17720# a_10616_17775# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X704 a_4681_16880# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X705 a_9736_15448# a_1692_17302# vssd1 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X706 vccd1 a_10092_5079# a_10004_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X707 vccd1 a_17820_3944# a_17732_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X708 vssd1 a_1772_6296# SDAC[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X709 a_26556_22760# a_26468_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X710 vccd1 a_13776_18100# a_14708_18100# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X711 a_24428_12919# a_24340_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X712 a_16120_23992# a_15156_23671# a_15916_23992# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X713 vssd1 a_1772_3160# SDAC[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X714 a_7190_18884# a_6358_19378# a_7022_18884# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X715 a_8455_13880# a_8335_13352# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X716 vccd1 a_11664_10704# a_11559_10304# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X717 vssd1 a_3564_20408# a_1772_20408# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X718 vssd1 a_13496_17337# a_11628_18056# vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X719 a_22372_25560# a_21204_25239# a_22168_25560# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X720 a_5836_22760# a_14649_21584# vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X721 a_12108_21664# a_15456_19368# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X722 a_12309_14180# a_12189_14136# a_11565_14136# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X723 vccd1 a_26668_16055# a_26580_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X724 vccd1 a_14895_24372# a_15351_24394# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X725 a_15025_21724# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X726 vccd1 a_26668_12919# a_26580_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X727 vccd1 a_16588_5079# a_16500_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X728 vccd1 a_24876_8215# a_24788_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X729 vccd1 a_19164_13352# a_19076_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X730 a_6396_3511# a_6308_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X731 a_13900_8215# a_13812_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X732 vccd1 a_14012_3944# a_13924_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X733 vssd1 a_24640_25940# DIGITAL_OUT[5] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X734 a_2444_24328# a_9920_20096# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X735 vccd1 a_14089_13744# a_13984_13884# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X736 vccd1 a_18604_11351# a_18516_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X737 a_13776_18100# a_11628_18056# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X738 a_20508_13352# a_20420_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X739 vssd1 a_16520_20128# a_6388_6390# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X740 a_5559_13016# a_5831_12568# a_4684_7564# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X741 a_20508_10216# a_20420_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X742 a_14708_18100# a_13776_18100# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X743 vssd1 a_2444_26249# COMP_CLK vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X744 vccd1 a_4481_24757# a_15324_25560# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X745 vssd1 a_13488_11000# a_3564_9432# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X746 vssd1 a_1772_9432# SDAC[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D15 a_1692_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X747 vccd1 a_22636_20759# a_22548_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X748 vccd1 a_13496_17337# a_11628_18056# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X749 a_14142_11850# a_13686_12404# a_13910_11850# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X750 vccd1 a_11548_3511# a_11460_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X751 vccd1 a_10876_5512# a_10788_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X752 a_5836_22760# a_14649_21584# vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X753 a_11856_25244# a_9332_25239# a_11544_25244# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X754 vccd1 a_11235_14136# a_9992_12846# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X755 a_27004_16488# a_26916_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X756 vccd1 a_13488_11000# a_3564_9432# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X757 vssd1 a_15456_19368# a_12108_21664# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X758 vssd1 a_15288_22021# a_14248_20686# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X759 a_21616_25560# a_21204_25239# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X760 vccd1 a_22076_21192# a_21988_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X761 a_7302_14180# a_6470_14674# a_7134_14180# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X762 vccd1 a_9196_5079# a_9108_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X763 a_28012_19191# a_27924_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X764 a_22636_9783# a_22548_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X765 a_9908_17016# a_5612_17317# vssd1 vssd1 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X766 a_28012_16055# a_27924_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X767 vccd1 a_23196_13352# a_23108_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X768 vccd1 a_23644_7080# a_23556_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X769 vccd1 a_22636_14487# a_22548_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D16 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X770 vccd1 a_3072_10564# a_5139_21292# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X771 vccd1 a_26556_19624# a_26468_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X772 a_7404_9006# a_1692_17302# a_8420_9176# vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X773 vccd1 a_22636_11351# a_22548_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X774 vccd1 a_7744_11088# a_7639_11459# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X775 vccd1 a_17372_7080# a_17284_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D17 vssd1 a_2140_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X776 a_16140_5079# a_16052_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X777 a_6215_21028# a_5759_20452# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X778 a_12650_11828# a_12026_11828# a_12502_12404# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X779 a_14895_24372# a_14271_24372# a_14747_24948# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X780 a_12189_14136# a_12581_14136# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X781 a_11212_6647# a_11124_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X782 vccd1 a_9920_20096# a_2444_24328# vccd1 pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X783 vccd1 a_25212_13352# a_25124_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X784 a_15804_11784# a_15716_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X785 a_10500_25560# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X786 a_24876_12919# a_24788_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X787 SDAC[6] a_1772_23544# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X788 a_3024_23292# a_2876_22848# a_2856_23292# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X789 vssd1 a_11076_24372# a_14271_22804# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X790 vccd1 a_3484_5512# a_3396_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X791 a_13364_12612# a_9444_19668# a_12581_14136# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X792 a_7337_25940# a_6607_25962# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X793 SDAC[5] a_1772_20408# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X794 a_3024_20156# a_2876_19712# a_2856_20156# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X795 vssd1 a_13832_15424# a_5612_17317# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X796 a_14403_24328# a_14068_23992# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X797 vccd1 a_10900_14964# a_1692_17302# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X798 a_2968_17317# a_3228_17317# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X799 vssd1 a_8156_17584# a_6328_17342# vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X800 a_27004_22327# a_26916_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X801 a_24092_19624# a_24004_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X802 SDAC[1] a_1772_6296# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X803 vccd1 a_2876_22848# a_2772_22892# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X804 a_11628_18056# a_13496_17337# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X805 a_27452_25896# a_27364_25940# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X806 a_17785_23632# a_17368_23676# a_18161_23676# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X807 SDAC[0] a_1772_3160# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X808 a_10716_22848# a_10408_22892# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X809 vssd1 a_23644_23291# a_23556_23335# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X810 a_20956_13352# a_20868_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X811 a_4152_12316# a_2352_11899# a_3212_11872# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X812 a_14708_18100# a_13776_18100# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X813 a_13564_5512# a_13476_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X814 a_20956_10216# a_20868_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X815 a_6630_18884# a_6154_19460# a_6358_19378# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X816 a_17372_18056# a_17284_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X817 a_10500_13016# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X818 COMP_CLK a_2444_26249# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X819 vccd1 a_23084_19191# a_22996_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X820 a_12543_14964# a_11919_14964# a_12375_14964# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X821 a_17372_14920# a_17284_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X822 vccd1 a_19500_17623# a_19412_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X823 vccd1 a_17932_12919# a_17844_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X824 vssd1 a_5836_22760# a_7628_20155# vssd1 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X825 vccd1 a_19276_8215# a_19188_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D18 vssd1 a_2444_24328# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X826 a_20620_9783# a_20532_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X827 a_11760_11828# a_10787_11829# vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X828 a_11548_13824# a_13496_15774# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X829 vccd1 a_2876_13440# a_2772_13484# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X830 vccd1 a_22748_3944# a_22660_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X831 vssd1 a_20652_22424# a_25648_25560# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D19 vssd1 a_1692_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X832 a_4760_12613# a_5020_12613# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X833 a_27452_16488# a_27364_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X834 a_4200_9180# a_3360_8763# a_3912_8780# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X835 vccd1 a_2876_10304# a_2772_10348# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X836 vssd1 a_15456_19368# a_12108_21664# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X837 vccd1 a_21404_19624# a_21316_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X838 a_12189_14136# a_12581_14136# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X839 a_9980_5512# a_9892_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X840 a_1772_9432# a_3564_9432# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X841 a_2568_22892# a_2016_22875# a_2364_22892# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X842 a_14232_21724# a_12020_21720# a_13292_21280# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X843 a_12085_16324# a_11965_15704# a_11341_15704# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X844 a_7758_10282# a_7302_10836# a_7526_10282# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X845 vccd1 a_7485_15496# a_7605_14964# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X846 vssd1 a_12413_11000# a_12533_11044# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X847 a_12444_3511# a_12356_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X848 a_17260_16055# a_17172_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X849 a_11076_24372# a_10372_24372# vccd1 vccd1 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X850 vccd1 a_16744_22042# a_10452_18840# vccd1 pfet_06v0 ad=0.458p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X851 a_14000_20856# a_13588_20535# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X852 vccd1 a_3324_16576# a_3220_16620# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X853 a_5880_12288# a_5860_14964# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X854 vssd1 a_1772_15704# SDAC[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X855 a_12085_15748# a_11965_15704# a_11341_15704# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X856 a_6172_5512# a_6084_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X857 vccd1 a_24540_24328# a_24452_24372# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X858 vccd1 a_18268_10216# a_18180_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X859 vccd1 a_4481_24757# a_7484_23992# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X860 a_8836_24372# a_8132_24372# vccd1 vccd1 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X861 a_7804_9831# a_7496_9880# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X862 a_6742_14180# a_6266_14756# a_6470_14674# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X863 a_2568_13484# a_2016_13467# a_2364_13484# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X864 vccd1 a_24092_16488# a_24004_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X865 vccd1 a_25660_13352# a_25572_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X866 vccd1 a_10764_6647# a_10676_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X867 a_17036_9783# a_16948_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X868 a_14872_25615# a_14471_25571# a_13815_25380# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X869 vccd1 a_23532_17623# a_23444_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X870 a_13116_7080# a_13028_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X871 a_2568_10348# a_2016_10331# a_2364_10348# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X872 a_10378_18884# a_4815_20408# a_10174_18884# vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X873 a_10296_25560# a_9332_25239# a_10092_25560# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X874 a_2276_22424# a_1828_22065# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X875 vssd1 a_4481_24757# a_12499_20152# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.217p ps=1.515u w=0.36u l=0.6u
X876 a_10472_14181# a_8617_15448# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X877 DIGITAL_OUT[0] a_9408_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X878 a_15916_23992# a_15816_23822# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X879 vccd1 a_3072_10564# a_10555_10216# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X880 a_24876_5079# a_24788_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X881 a_27452_22327# a_27364_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X882 vccd1 a_15244_5079# a_15156_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X883 vccd1 a_23532_8215# a_23444_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D20 a_2220_24686# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X884 a_2352_11899# a_1940_12312# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X885 a_18256_25560# a_17844_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X886 a_21292_19191# a_21204_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D21 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X887 a_21292_16055# a_21204_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X888 a_2016_22875# a_1604_23288# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X889 a_7829_8484# a_7709_7864# a_7085_7864# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X890 a_3999_21676# a_4233_23152# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X891 vccd1 a_19276_14487# a_19188_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X892 vssd1 a_18256_25560# DIGITAL_OUT[3] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X893 a_22300_16488# a_22212_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X894 a_27116_12919# a_27028_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X895 a_19164_3944# a_19076_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X896 a_7281_7142# a_2140_17302# a_7301_7608# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X897 vccd1 a_14460_3944# a_14372_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X898 vssd1 a_13776_18100# a_14708_18100# vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X899 a_20508_5512# a_20420_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X900 a_16140_8648# a_16052_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X901 vccd1 a_10372_24372# a_11076_24372# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X902 vccd1 a_8492_24328# a_8336_24372# vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
D22 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X903 a_8300_3511# a_8212_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X904 vccd1 a_2444_26249# COMP_CLK vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X905 a_16388_25940# a_15940_26471# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X906 a_20508_19624# a_20420_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X907 a_4233_15312# a_3816_15452# a_4609_15452# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X908 a_9900_13396# a_9444_13880# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X909 a_4464_12316# a_2352_11899# a_4152_12316# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X910 vccd1 a_10204_3511# a_10116_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X911 vccd1 a_6635_11000# a_6547_11045# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X912 vccd1 a_18156_16055# a_18068_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X913 a_11656_23292# a_9856_22875# a_10716_22848# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X914 vccd1 a_21852_19624# a_21764_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X915 vccd1 a_20060_14920# a_19972_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X916 a_19408_23992# a_19308_23544# vccd1 vccd1 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X917 vccd1 a_6154_19460# a_6590_19460# vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X918 a_2016_13467# a_1604_13880# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X919 vccd1 a_7804_9831# a_7700_9880# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X920 a_6983_11268# a_7639_11459# a_7535_11503# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X921 vccd1 a_20060_11784# a_19972_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X922 a_4609_18588# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X923 vccd1 a_9868_6647# a_9780_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X924 vccd1 a_16140_10216# a_16052_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X925 a_5895_21372# a_5795_21280# a_4771_21192# vccd1 pfet_06v0 ad=0.27805p pd=2.17u as=0.1079p ps=0.935u w=0.415u l=0.5u
D23 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X926 a_16924_3511# a_16836_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X927 vccd1 a_11996_3511# a_11908_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X928 a_12108_21664# a_15456_19368# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X929 vccd1 a_22300_7080# a_22212_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X930 vssd1 a_3072_10564# a_11043_10748# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X931 a_7123_11124# a_6983_11268# a_6635_11000# vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X932 vccd1 XRST a_7540_3249# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X933 a_8212_8693# a_1692_17302# a_7404_9006# vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X934 vccd1 a_1692_18885# a_1604_18929# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X935 vccd1 a_25324_23895# a_25236_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X936 a_10468_20152# a_7259_24800# a_9444_19668# vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X937 SDAC[6] a_1772_23544# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X938 vccd1 a_6271_22596# a_6727_22574# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X939 vccd1 a_25324_20759# a_25236_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X940 a_13116_3511# a_13028_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X941 vssd1 a_25648_25560# EOC vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X942 DIGITAL_OUT[4] a_21392_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X943 vssd1 a_12636_21976# a_12100_22020# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X944 vccd1 a_23980_17623# a_23892_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X945 a_13900_12568# a_10871_12268# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X946 vssd1 a_3999_21676# a_5647_22020# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X947 vccd1 a_2140_8648# a_2052_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X948 a_11412_21720# a_11292_21192# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X949 a_7205_8462# a_7085_7864# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X950 vccd1 a_2140_5512# a_2052_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X951 a_23644_8648# a_23556_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X952 a_5524_23288# a_5836_22760# a_3404_24812# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X953 vssd1 a_19648_21976# a_3564_25112# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X954 vccd1 a_22188_16055# a_22100_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X955 a_22372_25560# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X956 a_20280_24860# a_19352_24460# a_20112_24860# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X957 vssd1 a_6531_13789# a_6239_12568# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X958 a_19612_13352# a_19524_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X959 a_7628_20155# a_4815_20408# vssd1 vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X960 a_6499_21264# a_5795_21280# a_6915_21324# vccd1 pfet_06v0 ad=0.19315p pd=1.27u as=0.101p ps=0.905u w=0.505u l=0.5u
X961 vccd1 a_22188_12919# a_22100_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X962 vssd1 a_12413_9432# a_12533_9476# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X963 vccd1 a_25324_14487# a_25236_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X964 a_17372_8648# a_17284_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X965 a_19612_10216# a_19524_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X966 a_10787_11829# a_7988_19668# a_10599_11829# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X967 vccd1 a_19724_5079# a_19636_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X968 a_11660_6647# a_11572_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X969 a_7496_9880# a_6944_9880# a_7292_9880# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X970 vccd1 a_25324_11351# a_25236_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X971 a_11960_10348# a_11664_10704# a_10903_10216# vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X972 a_8645_10744# a_1692_17302# a_8437_10291# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X973 vssd1 a_3564_15704# a_1772_15704# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X974 a_2700_11916# a_2600_11872# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X975 vccd1 a_9308_3511# a_9220_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X976 vccd1 a_14124_11351# a_14036_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D24 vssd1 a_2444_24328# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X977 a_8009_22804# a_7279_22826# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X978 a_1916_22021# a_5836_22760# vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X979 vccd1 a_11965_15704# a_12085_16324# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
D25 vssd1 a_2444_24328# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X980 vccd1 a_11628_18056# a_9800_18056# vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X981 vccd1 a_20508_16488# a_20420_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X982 a_12579_24765# a_12909_24837# a_13029_24394# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
D26 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X983 a_12220_5512# a_12132_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X984 a_8492_11448# a_8040_11503# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X985 a_15064_25502# a_14576_25200# a_15324_25560# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X986 a_2096_24372# a_2220_24686# a_2116_24856# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X987 a_27564_12919# a_27476_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X988 a_17024_25940# a_16388_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X989 vccd1 a_22412_18056# a_22324_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X990 a_19276_5079# a_19188_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D27 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X991 a_7055_22804# a_6431_22804# a_6887_22804# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X992 vssd1 a_11965_15704# a_12085_15748# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X993 vccd1 a_2444_26249# COMP_CLK vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X994 a_3507_21237# a_2500_22020# a_3527_21720# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X995 a_20956_19624# a_20868_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X996 a_18716_5512# a_18628_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X997 a_26108_3944# a_26020_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X998 vccd1 a_21404_3944# a_21316_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X999 a_22524_21192# a_22436_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1000 vccd1 a_6328_17342# a_1692_10688# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1001 a_14348_6647# a_14260_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1002 vccd1 a_3564_25112# a_1772_25112# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1003 vssd1 a_1692_18528# a_1604_23288# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1004 a_5685_16533# a_4681_16880# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1005 a_11235_14136# a_11565_14136# a_11685_14734# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1006 a_23644_13352# a_23556_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1007 a_16812_11351# a_16724_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1008 a_8617_15448# a_8721_14920# a_8225_14965# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1009 vccd1 a_6172_9432# a_4965_14136# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X1010 vccd1 a_8300_8648# a_8437_10291# vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1011 vccd1 a_8454_21572# a_3703_18840# vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1012 a_23644_10216# a_23556_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1013 a_4828_3944# a_4740_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1014 a_11100_3511# a_11012_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1015 a_8076_5512# a_7988_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1016 vssd1 a_4041_24812# a_3972_24860# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X1017 vssd1 a_3072_10564# a_3024_15452# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1018 vccd1 a_25772_23895# a_25684_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1019 a_12308_22020# a_9076_15704# a_12308_22424# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1020 a_3192_12316# a_2352_11899# a_2904_11916# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1021 vccd1 a_22188_8215# a_22100_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1022 a_18171_20452# a_7225_22424# a_9263_20408# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1023 a_4069_11598# a_3949_11000# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1024 a_9856_22875# a_9444_23288# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1025 vccd1 a_25772_20759# a_25684_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1026 vccd1 a_3816_20156# a_4233_20016# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1027 vssd1 a_14403_24328# a_14271_24372# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
D28 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1028 a_9444_19668# a_5836_22760# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1029 vccd1 a_3564_15704# a_1772_15704# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1030 a_2052_25940# a_1604_26471# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1031 vccd1 a_13496_15774# a_11548_13824# vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1032 vccd1 a_3564_12568# a_1772_12568# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1033 a_4220_8736# a_3912_8780# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1034 vccd1 a_15064_12613# a_8300_8648# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1035 a_3360_8763# a_2948_9176# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1036 vssd1 a_1772_25112# SC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1037 a_19477_21236# a_19357_21768# a_18733_21701# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1038 a_3207_19288# a_3887_18840# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1039 a_7485_15496# a_1872_14602# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1040 a_19352_24460# a_18951_24416# a_18295_24328# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1041 vccd1 a_5573_11829# a_8225_14965# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1042 vccd1 a_1692_17302# a_8437_10291# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X1043 a_10204_22892# a_10104_22848# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1044 a_10759_21720# a_1916_17302# a_10575_21720# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1045 vccd1 a_25772_14487# a_25684_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1046 a_27900_3944# a_27812_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1047 a_6499_21264# a_5547_21551# a_6935_21724# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X1048 a_3024_18588# a_2876_18144# a_2856_18588# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1049 vssd1 a_1692_10688# a_2052_17016# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1050 vccd1 a_25772_11351# a_25684_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1051 a_23532_5079# a_23444_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1052 a_13564_7080# a_13476_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1053 a_17484_9783# a_17396_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1054 vccd1 a_14572_11351# a_14484_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D29 a_2444_24328# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1055 vssd1 a_2444_24328# a_13252_22804# vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1056 vssd1 a_6154_19460# a_6630_18884# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1057 vccd1 a_6440_18056# a_1692_18528# vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1058 a_15595_15448# a_9900_13396# a_8852_15704# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1059 vccd1 a_9900_24756# a_21684_22020# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1060 SDAC[5] a_1772_20408# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1061 vccd1 a_19164_19191# a_19076_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1062 vccd1 a_20956_16488# a_20868_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1063 a_17368_23676# a_15568_23992# a_16428_23943# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
D30 vssd1 COMP_OUT diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1064 a_14708_18100# a_13776_18100# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X1065 a_21068_18056# a_20980_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1066 a_24092_14920# a_24004_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1067 a_16700_5512# a_16612_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1068 vccd1 a_26220_17623# a_26132_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1069 a_10324_13396# a_9076_15704# a_10136_13396# vccd1 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X1070 vccd1 a_15692_5079# a_15604_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1071 vccd1 a_12108_6647# a_12020_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1072 a_3072_10564# a_9744_8392# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1073 vccd1 a_23980_8215# a_23892_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1074 a_7700_9880# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1075 vssd1 a_9800_18056# a_8156_17584# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1076 vccd1 a_22860_18056# a_22772_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D31 a_2444_24328# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1077 vssd1 a_19357_21768# a_19477_21812# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1078 a_13496_15774# a_14708_18100# vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1079 vssd1 a_17844_25560# a_18256_25560# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1080 a_26243_24765# a_26573_24837# a_26693_24394# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1081 a_18403_21629# a_18733_21701# a_18853_21811# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1082 a_22972_21192# a_22884_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1083 a_1892_14180# a_2220_14136# a_1872_14602# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1084 a_18828_6647# a_18740_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1085 vccd1 a_16388_25940# a_17024_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1086 vssd1 a_3564_6296# a_1772_6296# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1087 a_1892_11044# a_2220_11000# a_1872_11466# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1088 a_18984_22021# a_3999_21676# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1089 vccd1 a_19612_3944# a_19524_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1090 vccd1 a_20172_8215# a_20084_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1091 vssd1 a_3564_3160# a_1772_3160# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1092 a_20956_5512# a_20868_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1093 vccd1 a_8524_6647# a_8436_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1094 vccd1 a_18268_14920# a_18180_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1095 a_17036_14487# a_16948_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1096 vccd1 a_10652_3511# a_10564_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1097 a_11324_19624# a_11348_22065# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1098 vccd1 a_18268_11784# a_18180_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D32 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1099 a_2220_14136# a_4716_18840# a_4180_18884# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1100 a_1692_10688# a_6328_17342# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1101 vccd1 a_12860_21976# a_12736_22424# vccd1 pfet_06v0 ad=0.6588p pd=3.52u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1102 vccd1 a_26668_8215# a_26580_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1103 a_9076_15704# a_5019_20408# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1104 vccd1 a_1692_10688# a_2052_17016# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1105 vssd1 a_7709_7864# a_7829_7908# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1106 a_6915_21324# a_5895_21372# vccd1 vccd1 pfet_06v0 ad=0.101p pd=0.905u as=0.3975p ps=2.185u w=0.505u l=0.5u
X1107 a_6328_17342# a_8156_17584# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1108 vccd1 a_18716_13352# a_18628_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1109 a_21740_9783# a_21652_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1110 a_7055_11828# a_6431_11828# a_6907_12404# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1111 vccd1 a_20620_14487# a_20532_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1112 vccd1 a_13900_9783# a_13812_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1113 vccd1 a_11459_9432# a_10159_10700# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1114 vccd1 a_3072_10564# a_6635_11000# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X1115 a_12413_9432# a_8752_8648# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1116 a_14344_20156# a_13416_19756# a_14176_20156# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1117 vccd1 a_24540_19624# a_24452_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1118 a_15456_19368# a_14708_18100# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1119 vccd1 a_13900_6647# a_13812_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1120 a_10348_17016# a_8736_19363# a_10036_16532# vssd1 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1121 vccd1 a_13494_14136# a_1916_17302# vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1122 vccd1 a_27004_10216# a_26916_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1123 a_14475_22020# a_13999_22596# a_14223_22020# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1124 a_2568_15052# a_1604_15448# a_2364_15052# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1125 vssd1 a_8927_13836# a_8863_13880# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
D33 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1126 a_22300_8648# a_22212_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1127 a_10696_23292# a_9856_22875# a_10408_22892# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1128 a_13564_3511# a_13476_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1129 vssd1 a_7452_21280# a_7348_21324# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1130 vccd1 a_12668_5512# a_12580_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1131 a_27317_24948# a_27197_24904# a_26573_24837# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1132 vccd1 a_28012_23895# a_27924_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1133 vccd1 CLK a_13496_17337# vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1134 vccd1 a_28012_20759# a_27924_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1135 vssd1 a_9800_14181# a_2220_11000# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1136 a_26693_24947# a_26573_24837# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1137 a_9076_15704# a_5836_22760# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X1138 a_8624_14602# a_4348_7909# vccd1 vccd1 pfet_06v0 ad=0.4012p pd=1.85u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1139 a_24428_9783# a_24340_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1140 a_9479_10261# a_10159_10700# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1141 a_6736_23632# a_1692_18528# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1142 a_13048_16576# a_12560_16976# a_13308_16620# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1143 a_20508_7080# a_20420_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1144 vccd1 a_21628_21192# a_21540_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1145 a_19612_19624# a_19524_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1146 a_24428_17623# a_24340_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1147 a_6553_24373# a_5817_24800# vccd1 vccd1 pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1148 vccd1 a_4233_23152# a_4128_23292# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1149 vssd1 a_9800_18056# a_8156_17584# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1150 vccd1 a_9756_3511# a_9668_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1151 vssd1 a_3564_25112# a_1772_25112# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1152 a_8454_21572# a_8940_21590# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X1153 vssd1 a_14649_21584# a_14544_21724# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1154 vccd1 a_22748_13352# a_22660_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1155 SDAC[1] a_1772_6296# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1156 vccd1 a_19164_7080# a_19076_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1157 vssd1 a_11787_20027# a_9920_20096# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1158 vccd1 a_7597_15704# a_7717_16324# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1159 SDAC[0] a_1772_3160# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1160 a_19164_11784# a_19076_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1161 vssd1 a_21392_25940# DIGITAL_OUT[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1162 a_8435_13397# a_8519_13836# a_8455_13880# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1163 a_3619_11000# a_3949_11000# a_4069_11598# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1164 a_20652_22424# a_20196_22112# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1165 vccd1 a_28012_14487# a_27924_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1166 vccd1 a_22636_5079# a_22548_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1167 vccd1 a_16388_25940# a_17024_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1168 a_9744_8392# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X1169 vccd1 a_28012_11351# a_27924_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1170 vccd1 a_3703_18840# a_5559_11448# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
D34 CLK vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1171 a_20060_3944# a_19972_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1172 a_5500_13352# a_5412_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1173 vssd1 a_7597_15704# a_7717_15748# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1174 a_20508_14920# a_20420_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1175 vccd1 a_5276_5512# a_5188_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1176 a_19500_20759# a_19412_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1177 vccd1 a_18380_8215# a_18292_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1178 a_24640_25940# a_24004_22804# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1179 a_17484_14487# a_17396_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1180 vccd1 a_4233_13744# a_4128_13884# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1181 a_8153_25200# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1182 a_23725_24904# a_20260_23588# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1183 vccd1 a_4233_10608# a_4128_10748# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1184 vssd1 a_5084_25560# a_13216_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1185 a_1996_11000# a_10584_22042# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X1186 a_5057_17020# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1187 a_26556_3944# a_26468_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1188 vccd1 a_21852_3944# a_21764_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1189 a_14796_6647# a_14708_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1190 a_1692_10688# a_6328_17342# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1191 a_22188_5079# a_22100_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1192 vssd1 a_1692_17302# a_9540_12268# vssd1 nfet_06v0 ad=0.104p pd=0.92u as=0.14p ps=1.1u w=0.4u l=0.6u
X1193 vccd1 a_15456_19368# a_12108_21664# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1194 vccd1 a_1692_10688# a_1940_12312# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1195 a_9420_6647# a_9332_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1196 a_23644_19624# a_23556_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1197 vssd1 a_3564_12568# a_1772_12568# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1198 a_25212_21192# a_25124_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1199 a_11628_18056# a_13496_17337# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1200 vccd1 a_8524_5512# a_8436_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1201 a_15356_5512# a_15268_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1202 a_12340_18884# a_10555_21267# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1203 a_3072_10564# a_9744_8392# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X1204 a_4752_7864# a_4716_18840# vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X1205 a_19500_11351# a_19412_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1206 a_23196_11784# a_23108_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D35 a_5940_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1207 vccd1 a_27452_10216# a_27364_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D36 XRST vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1208 a_23728_25244# a_21616_25560# a_23416_25244# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1209 vccd1 a_22636_19191# a_22548_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1210 a_4693_17316# a_4573_17272# a_3949_17272# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1211 vccd1 a_19612_16488# a_19524_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1212 a_8841_20152# a_8144_19288# a_7932_20453# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1213 a_6719_16532# a_6095_16532# a_6551_16532# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
D37 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1214 vccd1 a_22157_23336# a_22277_22804# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1215 a_3703_18840# a_8454_21572# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1216 vssd1 a_3507_21237# a_5423_19668# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1217 a_12220_7080# a_12132_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1218 vccd1 a_13900_8648# a_13812_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1219 a_16140_9783# a_16052_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1220 a_21964_25560# a_21864_25390# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
D38 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1221 a_23532_20759# a_23444_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1222 vccd1 a_18268_3944# a_18180_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1223 a_7225_22424# a_6495_22020# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X1224 a_25212_11784# a_25124_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1225 a_11544_25244# a_9744_25560# a_10604_25511# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1226 a_19357_18632# a_5020_15796# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1227 a_11628_18056# a_13496_17337# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1228 vccd1 a_20620_5079# a_20532_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1229 a_24876_17623# a_24788_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1230 a_23084_12919# a_22996_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1231 EOC a_25648_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1232 a_18716_7080# a_18628_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1233 a_23980_5079# a_23892_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1234 a_5860_14964# a_5412_15495# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1235 a_14348_8215# a_14260_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1236 a_16812_16055# a_16724_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D39 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1237 vssd1 a_21392_25940# DIGITAL_OUT[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1238 vssd1 a_9900_24756# a_18996_23588# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1239 vccd1 a_24316_22327# a_24228_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1240 a_3228_17317# a_1804_21723# a_3207_19288# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1241 a_23532_14487# a_23444_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1242 a_16520_20128# COMP_OUT vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1243 a_8352_23676# a_6736_23632# a_7224_23934# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1244 a_22277_23380# a_22157_23336# a_21533_23269# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1245 a_10740_16532# a_10036_16532# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1246 a_23532_11351# a_23444_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1247 a_24540_3944# a_24452_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1248 vccd1 a_26108_7080# a_26020_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1249 vccd1 a_17260_11351# a_17172_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1250 a_8433_20152# a_7337_20856# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1251 vccd1 a_12556_6647# a_12468_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1252 a_8868_14609# a_8519_13836# a_8624_14602# vccd1 pfet_06v0 ad=0.58035p pd=2.155u as=0.4012p ps=1.85u w=1.095u l=0.5u
X1253 a_20172_5079# a_20084_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1254 a_19556_23992# a_18996_23588# a_19428_23588# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X1255 a_11939_17020# a_11799_16488# a_11451_16488# vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X1256 a_20956_14920# a_20868_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1257 vssd1 a_1772_6296# SDAC[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1258 vccd1 a_23644_16488# a_23556_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1259 vssd1 a_1772_3160# SDAC[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1260 vccd1 a_10192_8692# a_4481_24757# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1261 a_10820_20452# a_9920_20096# a_10616_20452# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1262 a_2788_19288# a_1996_11000# a_2544_19306# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X1263 a_14727_24372# a_14271_24372# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1264 a_4751_20452# a_4631_20408# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1265 a_26668_5079# a_26580_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1266 vccd1 a_17036_5079# a_16948_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1267 a_12780_21324# a_11392_21236# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1268 vccd1 a_21292_20759# a_21204_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1269 a_9444_19668# a_9532_19624# vccd1 vccd1 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1270 vccd1 a_15456_19368# a_12108_21664# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1271 vccd1 a_25324_8215# a_25236_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1272 a_13497_14964# a_12767_14986# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1273 vccd1 a_22300_10216# a_22212_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1274 a_16408_23676# a_15568_23992# a_16120_23992# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1275 vccd1 a_2876_18144# a_2772_18188# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1276 a_5559_13016# a_6239_12568# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1277 vccd1 a_8972_6647# a_8884_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1278 a_25660_21192# a_25572_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1279 a_5160_9180# a_3360_8763# a_4220_8736# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1280 vssd1 a_14428_23544# a_14380_23588# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X1281 vccd1 a_17368_23676# a_17785_23632# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1282 vssd1 a_14652_12605# a_14350_13016# vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1283 vccd1 a_15804_3511# a_15716_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1284 a_5880_12288# a_5860_14964# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1285 vccd1 a_18256_25560# DIGITAL_OUT[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1286 vssd1 a_4233_13744# a_4128_13884# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1287 a_5237_13397# a_4233_13744# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1288 a_5577_9040# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
D40 a_2444_24328# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1289 vssd1 a_1916_17302# a_1812_17353# vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1290 a_5237_10261# a_4233_10608# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1291 vccd1 a_16252_3944# a_16164_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1292 vssd1 a_4233_10608# a_4128_10748# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1293 vccd1 a_18828_14487# a_18740_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1294 vccd1 a_21292_14487# a_21204_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1295 vccd1 a_21292_11351# a_21204_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1296 vssd1 a_13776_18100# a_14708_18100# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1297 vccd1 a_11324_5512# a_11236_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1298 vccd1 a_27900_7080# a_27812_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1299 COMP_CLK a_2444_26249# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1300 a_26668_23895# a_26580_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1301 vccd1 a_5076_23992# a_12132_19288# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X1302 a_23980_20759# a_23892_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1303 a_16700_7080# a_16612_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1304 a_9444_19668# a_9920_20096# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1305 vccd1 a_17708_16055# a_17620_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1306 a_14652_12605# a_14089_13744# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1307 a_25660_11784# a_25572_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1308 vssd1 a_17632_21976# a_5019_20408# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1309 a_2568_18188# a_2016_18171# a_2364_18188# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1310 vssd1 a_5237_18101# a_5530_18884# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1311 a_11628_18056# a_13496_17337# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D41 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1312 vccd1 a_20172_12919# a_20084_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1313 a_18716_3511# a_18628_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1314 a_25648_25560# a_20652_22424# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1315 vccd1 a_4731_20872# a_6060_23118# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1316 a_9560_20452# a_9920_20096# a_11248_20452# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1317 a_18828_8215# a_18740_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1318 a_12108_21664# a_15456_19368# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1319 SDAC[4] a_1772_15704# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1320 vccd1 a_11459_11000# a_11279_12268# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1321 vccd1 a_24764_22327# a_24676_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1322 vssd1 a_12189_14136# a_12309_14180# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1323 a_23980_14487# a_23892_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1324 a_4828_5079# a_4740_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1325 a_8076_6647# a_7988_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1326 vssd1 a_17859_24373# a_19748_26471# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1327 a_20956_7080# a_20868_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1328 a_24876_9783# a_24788_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1329 vccd1 a_11451_16488# a_5020_15796# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1330 a_23980_11351# a_23892_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1331 vccd1 a_9123_17317# a_10900_14964# vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1332 vccd1 a_1772_23544# SDAC[6] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1333 vccd1 a_4152_12316# a_4569_12176# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
D42 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1334 DIGITAL_OUT[4] a_21392_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1335 a_5940_6390# a_12262_23544# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1336 vccd1 a_1772_20408# SDAC[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1337 a_11459_9432# a_11789_9432# a_11909_10030# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1338 a_14736_20156# a_13015_19712# a_13608_19712# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1339 a_9444_19668# a_7259_24800# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1340 a_18380_5079# a_18292_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1341 vccd1 a_24316_21192# a_24228_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1342 a_27116_17623# a_27028_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1343 a_13815_25380# a_14576_25200# a_14367_25615# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X1344 a_17820_5512# a_17732_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1345 a_19164_8648# a_19076_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1346 SC a_1772_25112# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1347 a_25212_3944# a_25124_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1348 a_2444_24328# a_9920_20096# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X1349 a_13452_6647# a_13364_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D43 vssd1 a_2220_24686# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1350 vccd1 a_13686_12404# a_14142_11850# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1351 a_14747_23380# a_14271_22804# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1352 vccd1 a_27004_14920# a_26916_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1353 vccd1 a_6396_3511# a_6308_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1354 SDAC[1] a_1772_6296# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1355 a_10092_25560# a_8836_24372# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1356 a_3016_16620# a_2464_16603# a_2812_16620# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1357 SDAC[0] a_1772_3160# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1358 vssd1 a_2444_24328# a_20859_26424# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1359 a_18295_24328# a_18951_24416# a_18847_24460# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1360 vssd1 a_5237_13397# a_5642_14180# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1361 vccd1 a_27004_11784# a_26916_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1362 vccd1 a_20060_19624# a_19972_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1363 a_27197_24904# a_23644_23291# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1364 vssd1 a_14068_23992# a_14403_24328# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1365 a_3932_3944# a_3844_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1366 a_14012_5512# a_13924_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1367 a_7180_5512# a_7092_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1368 a_4233_18448# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1369 vccd1 a_21292_8215# a_21204_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1370 vssd1 a_1692_10688# a_1940_12312# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1371 a_13868_19756# a_13416_19756# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X1372 a_10472_14181# a_8617_15448# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
D44 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1373 a_13955_25236# a_13815_25380# a_13467_25112# vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X1374 SDAC[4] a_1772_15704# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1375 a_6983_11268# a_7744_11088# a_7535_11503# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X1376 SDAC[3] a_1772_12568# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1377 vccd1 a_15804_5512# a_15716_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1378 vccd1 a_3507_21237# a_5423_19668# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1379 a_23196_3944# a_23108_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1380 a_7643_12612# a_7167_13188# a_7391_12612# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1381 a_4088_7909# a_4348_7909# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1382 vccd1 a_10192_8692# a_4481_24757# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1383 vccd1 a_3564_25112# a_1772_25112# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1384 vccd1 a_11787_20027# a_9920_20096# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1385 vccd1 a_8132_24372# a_8836_24372# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1386 vssd1 a_1692_18528# a_2724_24856# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1387 a_10716_22848# a_10408_22892# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1388 a_25648_25560# a_20652_22424# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1389 vccd1 a_5612_17317# a_5524_17361# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1390 a_23416_25244# a_21616_25560# a_22476_25511# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1391 vccd1 a_13496_17337# a_11628_18056# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1392 vccd1 a_25324_19191# a_25236_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1393 vssd1 a_6531_15357# a_2712_16576# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1394 a_6553_24373# a_5817_24800# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1395 a_7485_15496# a_1872_14602# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1396 a_19612_14920# a_19524_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D45 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1397 a_2700_11916# a_2600_11872# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
D46 a_2140_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1398 vccd1 a_17221_20453# a_20196_22112# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1399 a_3816_23292# a_1604_23288# a_2876_22848# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1400 a_6123_22020# a_5647_22020# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1401 vccd1 a_20060_7080# a_19972_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1402 a_26220_20759# a_26132_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1403 vccd1 a_3564_15704# a_1772_15704# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1404 vccd1 a_11212_6647# a_11124_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1405 a_10192_8692# a_7988_3608# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1406 a_11451_16488# a_11799_16488# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X1407 vccd1 a_13496_15774# a_11548_13824# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1408 a_14796_8215# a_14708_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D47 a_2220_24686# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1409 vccd1 a_3564_12568# a_1772_12568# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1410 a_4481_24757# a_10192_8692# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1411 a_11628_18056# a_13496_17337# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1412 a_12533_11620# a_12413_11000# a_11789_11000# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1413 DIGITAL_OUT[5] a_24640_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1414 a_27564_17623# a_27476_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1415 vssd1 a_10676_16152# a_11919_14964# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1416 vccd1 a_13216_25940# DIGITAL_OUT[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1417 a_7195_17107# a_6719_16532# a_6943_16554# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1418 vccd1 a_26556_7080# a_26468_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1419 vccd1 a_21392_25940# DIGITAL_OUT[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1420 a_17932_6647# a_17844_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1421 a_19276_9783# a_19188_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1422 a_4771_21192# a_5795_21280# a_5139_21292# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.2898p ps=2.33u w=0.36u l=0.6u
X1423 a_25324_5079# a_25236_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1424 a_15356_7080# a_15268_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1425 vccd1 a_27004_22327# a_26916_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D48 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1426 a_19500_16055# a_19412_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1427 vccd1 a_27452_14920# a_27364_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1428 vssd1 a_1772_6296# SDAC[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1429 vssd1 a_1692_18528# a_9332_25239# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1430 a_26220_14487# a_26132_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1431 a_10584_25244# a_9744_25560# a_10296_25560# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1432 vssd1 a_1772_3160# SDAC[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1433 a_6755_7864# a_7085_7864# a_7205_7908# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1434 a_26108_8648# a_26020_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1435 vccd1 a_27452_11784# a_27364_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1436 a_3816_13884# a_1604_13880# a_2876_13440# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1437 a_26220_11351# a_26132_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1438 vccd1 a_16252_11784# a_16164_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1439 vssd1 a_9408_25940# DIGITAL_OUT[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1440 a_3816_10748# a_1604_10744# a_2876_10304# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1441 a_15020_11351# a_14932_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1442 vccd1 a_18716_19191# a_18628_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1443 a_14465_13884# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1444 vccd1 a_7302_10836# a_7758_10282# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1445 a_7932_20453# a_8144_19288# a_8225_19669# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1446 vccd1 a_17484_5079# a_17396_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1447 a_2340_24372# a_2220_24686# a_2096_24372# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X1448 a_23644_14920# a_23556_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1449 vccd1 a_27900_13352# a_27812_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1450 vccd1 a_25772_8215# a_25684_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1451 a_9056_9564# a_6532_9559# a_8744_9564# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1452 vssd1 a_13608_19712# a_13416_19756# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1453 vccd1 a_4672_12657# a_4836_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
D49 a_6388_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1454 vssd1 a_4233_23152# a_4128_23292# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
D50 vssd1 CLK diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1455 a_14068_23992# a_9900_24756# a_13920_23992# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X1456 vssd1 a_17585_20856# a_18171_20452# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1457 a_5237_19669# a_4233_20016# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1458 vccd1 a_25212_18056# a_25124_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1459 a_11548_13824# a_13496_15774# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1460 vssd1 a_4233_20016# a_4128_20156# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1461 a_22748_5512# a_22660_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1462 vccd1 a_3703_18840# a_3319_21237# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1463 a_20396_17623# a_20308_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1464 a_8841_15448# a_8721_14920# a_8617_15448# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1465 a_9900_24756# a_13252_22804# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X1466 a_23532_19191# a_23444_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1467 vssd1 a_17024_25940# DIGITAL_OUT[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1468 a_23532_16055# a_23444_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1469 vccd1 a_12444_3511# a_12356_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1470 vccd1 a_11772_5512# a_11684_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1471 a_20508_19191# a_20420_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1472 vssd1 a_1772_23544# SDAC[6] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1473 vccd1 a_7337_20856# a_8225_19669# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1474 vssd1 a_6388_6390# a_2220_24686# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1475 a_3136_24443# a_2724_24856# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1476 a_5940_6390# a_12262_23544# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1477 a_7001_19668# a_6271_19690# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X1478 vccd1 a_25772_19191# a_25684_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1479 vccd1 a_18403_18493# a_16773_18528# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1480 a_27900_8648# a_27812_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1481 a_15244_10216# a_15156_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D51 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1482 a_23532_9783# a_23444_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1483 a_1692_18528# a_6440_18056# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1484 a_2588_3944# a_2500_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1485 vccd1 a_4481_24757# a_13467_25112# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X1486 a_13940_23588# a_13820_23544# vssd1 vssd1 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1487 vccd1 a_24540_7080# a_24452_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1488 SC a_1772_25112# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1489 a_6115_23668# a_5975_23812# a_5627_23544# vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
D52 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1490 a_21628_3511# a_21540_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1491 a_11628_18056# a_13496_17337# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1492 vssd1 a_1916_17302# a_15595_15448# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1493 vccd1 a_22300_14920# a_22212_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1494 a_10604_25511# a_10296_25560# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1495 vccd1 a_7259_24800# a_2444_24328# vccd1 pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1496 DIGITAL_OUT[5] a_24640_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1497 a_3507_21237# a_2164_21236# a_3319_21237# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1498 a_10740_16532# a_10036_16532# vccd1 vccd1 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1499 a_8433_15448# a_5573_11829# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1500 a_15356_3511# a_15268_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1501 vccd1 a_22300_11784# a_22212_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1502 vccd1 a_13216_25940# DIGITAL_OUT[1] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1503 a_3108_11916# a_1940_12312# a_2904_11916# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1504 vccd1 a_21740_5079# a_21652_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1505 vccd1 a_21392_25940# DIGITAL_OUT[4] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1506 a_8121_13016# a_7391_12612# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1507 a_10036_16532# a_8736_19363# a_9888_16532# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X1508 a_18295_24328# a_19056_24816# a_18847_24460# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X1509 vccd1 a_27452_22327# a_27364_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1510 a_21180_21192# a_21092_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1511 a_11461_16302# a_11341_15704# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1512 vccd1 a_4380_5512# a_4292_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1513 vssd1 a_9408_25940# DIGITAL_OUT[0] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1514 a_25660_3944# a_25572_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1515 a_21292_5079# a_21204_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1516 a_24316_22760# a_24228_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1517 a_1772_6296# a_3564_6296# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1518 vssd1 a_2052_25940# a_9408_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1519 SDAC[3] a_1772_12568# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1520 a_1772_3160# a_3564_3160# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1521 vccd1 a_27004_21192# a_26916_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1522 vssd1 a_13496_17337# a_11628_18056# vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1523 a_11965_15704# a_9123_17317# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1524 vccd1 a_24428_5079# a_24340_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1525 vccd1 a_9161_9520# a_9056_9564# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1526 vccd1 a_24428_16055# a_24340_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1527 vccd1 a_8300_3511# a_8212_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1528 a_14460_5512# a_14372_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1529 a_11455_10348# a_10555_10216# vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1530 a_18716_11784# a_18628_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1531 a_2116_24856# a_2444_24328# a_2096_24372# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1532 vccd1 a_7259_24800# a_5612_23118# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1533 vccd1 a_24428_12919# a_24340_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1534 vccd1 a_25660_18056# a_25572_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1535 vccd1 a_4815_20408# a_3004_21664# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1536 a_16588_12919# a_16500_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1537 vccd1 a_10732_24328# a_15940_26471# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1538 vssd1 a_14708_18100# a_13496_15774# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1539 a_3728_24460# a_3136_24443# a_3524_24460# vccd1 pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1540 a_23980_19191# a_23892_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1541 a_11965_15704# a_9123_17317# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1542 a_5817_24800# a_4913_24860# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X1543 a_23980_16055# a_23892_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1544 vccd1 a_16924_3511# a_16836_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1545 vccd1 a_23644_3944# a_23556_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1546 a_16588_6647# a_16500_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1547 a_7134_14180# a_6470_14674# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1548 a_14000_20856# a_13588_20535# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1549 vccd1 a_17372_3944# a_17284_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1550 DIGITAL_OUT[2] a_17024_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1551 a_15692_10216# a_15604_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1552 a_1692_18528# a_6440_18056# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1553 a_2876_15008# a_2568_15052# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1554 vccd1 a_13116_3511# a_13028_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1555 a_4385_24860# a_3728_24460# vssd1 vssd1 nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1556 a_17820_7080# a_17732_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1557 a_12736_22424# a_12636_21976# a_12308_22020# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1558 a_18984_22021# a_3999_21676# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1559 vssd1 a_11628_18056# a_9800_18056# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1560 a_13452_8215# a_13364_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1561 a_5137_24860# a_3136_24443# a_4913_24860# vccd1 pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X1562 a_22748_11784# a_22660_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1563 vccd1 a_4716_25204# a_4628_25248# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1564 a_14747_24948# a_14271_24372# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1565 a_5975_23812# a_6631_24003# a_6527_24047# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1566 a_1812_17720# a_1692_17302# vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1567 vccd1 a_6047_19668# a_6503_19690# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1568 a_8156_17584# a_9800_18056# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1569 vccd1 a_25212_7080# a_25124_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1570 a_19164_16488# a_19076_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D53 a_1804_21723# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1571 vccd1 a_11660_6647# a_11572_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1572 a_14012_7080# a_13924_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1573 vccd1 a_28012_19191# a_27924_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D54 vssd1 a_6388_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1574 a_18435_24860# a_18295_24328# a_17947_24328# vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X1575 a_20060_8648# a_19972_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1576 a_10040_20152# a_9920_20096# a_9846_20152# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X1577 a_7348_21324# a_5795_21280# a_6499_21264# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1578 a_5620_18584# a_4672_12657# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1579 a_2464_16603# a_2052_17016# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1580 vccd1 a_14708_18100# a_13496_15774# vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X1581 vccd1 a_3932_7080# a_3844_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1582 a_1692_26427# a_8153_25200# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1583 a_7988_19668# a_7540_20199# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1584 a_25772_5079# a_25684_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1585 DIGITAL_OUT[3] a_18256_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1586 vccd1 a_4233_18448# a_4128_18588# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1587 a_13496_17337# CLK vccd1 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.428p ps=2.02u w=0.82u l=0.5u
X1588 a_22636_12919# a_22548_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1589 vccd1 a_16140_5079# a_16052_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1590 vssd1 a_2052_25940# a_9408_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1591 a_26556_8648# a_26468_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1592 vccd1 a_27452_21192# a_27364_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1593 a_8736_19363# a_10452_18840# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X1594 vccd1 a_7709_7864# a_7829_8484# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1595 vssd1 a_1772_20408# SDAC[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1596 a_5020_12613# a_2140_17302# a_15120_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1597 a_22188_9783# a_22100_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1598 vccd1 a_9540_12268# a_4492_18840# vccd1 pfet_06v0 ad=0.389p pd=2.02u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1599 vccd1 a_24876_16055# a_24788_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1600 a_3360_12316# a_3212_11872# a_3192_12316# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1601 vccd1 a_24876_12919# a_24788_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1602 vccd1 a_14348_9783# a_14260_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1603 a_14756_20856# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1604 vccd1 a_17372_13352# a_17284_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1605 vccd1 a_14348_6647# a_14260_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1606 vccd1 a_23196_7080# a_23108_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1607 a_14872_25615# a_14576_25200# a_13815_25380# vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1608 a_12581_14136# a_9444_19668# a_13572_13016# vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1609 a_8156_17584# a_9800_18056# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1610 vssd1 a_3564_6296# a_1772_6296# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1611 a_3708_8780# a_3608_8736# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1612 vssd1 a_24004_22804# a_24640_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1613 a_13077_22805# a_12073_23152# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1614 a_19357_21768# a_17221_20453# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1615 vccd1 a_16812_11351# a_16724_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1616 a_7452_21280# a_5940_6390# a_8583_20856# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1617 vssd1 a_14708_18100# a_13496_15774# vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1618 vssd1 a_3564_3160# a_1772_3160# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1619 a_21404_5512# a_21316_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1620 DIGITAL_OUT[1] a_13216_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1621 a_22244_22424# a_9900_24756# a_22096_22424# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X1622 vccd1 a_2588_8215# a_2500_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1623 a_2892_18840# a_5237_19669# a_12340_18884# vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1624 a_23196_16488# a_23108_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1625 a_15848_20128# a_5237_19669# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1626 vccd1 a_11100_3511# a_11012_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1627 vccd1 a_19357_21768# a_19477_21236# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1628 vssd1 a_6440_18056# a_1692_18528# vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1629 a_23308_18056# a_23220_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1630 a_12579_24765# a_12909_24837# a_13029_24947# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1631 a_9295_22596# a_8671_22020# a_9147_22020# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1632 a_7605_14964# a_7485_15496# a_6861_15429# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1633 a_12533_11044# a_12413_11000# a_11789_11000# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1634 a_8736_19363# a_4815_20408# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1635 a_14089_13744# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1636 vccd1 a_27116_8215# a_27028_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1637 a_9263_20408# a_7225_22424# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1638 a_1772_12568# a_3564_12568# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1639 vssd1 a_10192_8692# a_4481_24757# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1640 vccd1 a_5160_9180# a_5577_9040# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1641 a_17820_3511# a_17732_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1642 vssd1 a_2164_21236# a_8841_20152# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1643 a_12158_11784# a_11961_12656# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1644 a_8040_11503# a_7744_11088# a_6983_11268# vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1645 vccd1 a_1692_18528# a_2724_24856# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1646 a_25212_16488# a_25124_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1647 vssd1 a_6328_17342# a_1692_10688# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1648 vccd1 a_5940_6390# a_2444_18840# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1649 vccd1 a_6531_15357# a_2712_16576# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1650 a_17932_8215# a_17844_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1651 vssd1 a_13467_25112# a_10732_24328# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1652 a_23084_17623# a_22996_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1653 a_5132_7564# a_4964_9880# a_5559_11448# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1654 vccd1 a_1692_26427# a_1604_26471# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1655 a_26220_19191# a_26132_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1656 a_3932_5079# a_3844_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1657 vssd1 a_3072_10564# a_9699_17396# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X1658 a_26220_16055# a_26132_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D55 a_6388_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1659 a_23980_9783# a_23892_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1660 a_10104_22848# a_5612_23118# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1661 a_14012_3511# a_13924_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1662 vccd1 a_13116_5512# a_13028_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1663 vssd1 a_5577_9040# a_5472_9180# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1664 a_9800_18056# a_11628_18056# vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1665 a_6755_7864# a_7085_7864# a_7205_8462# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1666 a_26108_13352# a_26020_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1667 a_2856_15452# a_2016_15035# a_2568_15052# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1668 a_26108_10216# a_26020_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1669 a_24540_8648# a_24452_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D56 vssd1 a_2444_24328# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1670 a_4752_15704# a_5020_15796# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X1671 a_8972_16177# a_8852_15704# vccd1 vccd1 pfet_06v0 ad=0.2847p pd=1.615u as=0.5913p ps=3.27u w=1.095u l=0.5u
X1672 a_20172_9783# a_20084_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1673 vssd1 a_14649_21584# a_5836_22760# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1674 vssd1 XRST a_7540_3249# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1675 a_13496_17337# CLK vccd1 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1676 vssd1 a_6635_11000# a_6547_11045# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1677 a_7093_16302# a_6973_15704# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1678 vccd1 a_9532_5512# a_9444_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1679 SDAC[1] a_1772_6296# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1680 a_10604_25511# a_10296_25560# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1681 vccd1 a_24509_23544# a_24629_24164# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1682 vssd1 a_1772_20408# SDAC[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1683 SDAC[0] a_1772_3160# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1684 a_26668_9783# a_26580_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1685 a_22748_7080# a_22660_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1686 vccd1 a_18828_9783# a_18740_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1687 a_4935_20452# a_4815_20408# a_4751_20452# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1688 a_19612_19191# a_19524_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1689 a_9532_19624# a_1692_17302# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X1690 vccd1 a_25648_25560# EOC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1691 a_25212_22327# a_25124_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1692 vccd1 a_2220_14136# a_2116_14584# vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1693 vccd1 a_18828_6647# a_18740_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1694 a_8156_17584# a_9800_18056# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1695 a_11628_18056# a_13496_17337# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1696 vssd1 a_24640_25940# DIGITAL_OUT[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1697 vccd1 a_2220_11000# a_2116_11448# vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1698 vccd1 a_1772_23544# SDAC[6] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1699 vssd1 a_24509_23544# a_24629_23588# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1700 DIGITAL_OUT[1] a_13216_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1701 DIGITAL_OUT[4] a_21392_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1702 a_14953_22424# a_14223_22020# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1703 a_5237_18101# a_4233_18448# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1704 vssd1 a_13900_12568# a_13364_12612# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
D57 vssd1 a_5940_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1705 vccd1 a_1772_20408# SDAC[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1706 vssd1 a_4233_18448# a_4128_18588# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1707 vccd1 a_24876_5079# a_24788_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1708 a_4716_18840# a_4233_15312# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1709 a_19612_5512# a_19524_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1710 a_7224_23934# a_6631_24003# a_7960_23676# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1711 a_23756_18056# a_23668_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1712 vccd1 a_17036_14487# a_16948_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1713 a_27004_3944# a_26916_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1714 vssd1 a_13999_22596# a_14475_22020# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X1715 vccd1 a_21292_19191# a_21204_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1716 vccd1 a_22300_3944# a_22212_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1717 a_15244_6647# a_15156_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1718 a_27004_22760# a_26916_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1719 vccd1 a_14348_8648# a_14260_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1720 a_10864_23292# a_10716_22848# a_10696_23292# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1721 vssd1 a_2444_24328# a_9659_9176# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1722 vssd1 a_11459_9432# a_10159_10700# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1723 a_7597_15704# a_4716_18840# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1724 vssd1 a_27197_24904# a_27317_24948# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1725 vccd1 a_27116_16055# a_27028_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1726 vccd1 a_11961_25200# a_11856_25244# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1727 a_9751_22574# a_9295_22596# a_9519_22020# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X1728 a_25660_16488# a_25572_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1729 vccd1 a_27116_12919# a_27028_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1730 a_5724_3944# a_5636_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1731 vccd1 a_2588_7080# a_2500_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1732 vssd1 a_4684_7564# a_2600_11872# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1733 a_26243_24765# a_26573_24837# a_26693_24947# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1734 vssd1 a_6328_17342# a_1692_10688# vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1735 a_6727_22574# a_6271_22596# a_6495_22020# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X1736 a_19276_12919# a_19188_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1737 a_3072_10564# a_9744_8392# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1738 a_9540_12268# a_9532_13685# vssd1 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.104p ps=0.92u w=0.4u l=0.6u
X1739 vccd1 a_23084_8215# a_22996_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1740 a_13776_18100# a_11628_18056# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1741 a_6719_16532# a_6095_16532# a_6571_17108# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1742 a_10296_25560# a_9744_25560# a_10092_25560# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1743 a_18853_18122# a_18733_18565# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1744 a_4069_14180# a_3949_14136# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1745 a_3212_11872# a_2904_11916# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1746 vssd1 a_2444_26249# COMP_CLK vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1747 a_3108_11916# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1748 a_7205_7908# a_7085_7864# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1749 vssd1 a_13496_15774# a_11548_13824# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1750 a_19724_14487# a_19636_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1751 a_14350_13016# a_2140_17302# vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1752 vccd1 a_13564_3511# a_13476_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1753 a_4069_11044# a_3949_11000# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1754 vssd1 a_3619_14136# a_2264_13440# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1755 a_26556_13352# a_26468_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1756 a_8247_13397# a_8927_13836# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1757 a_26556_10216# a_26468_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1758 vssd1 a_3619_11000# a_2264_10304# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1759 vccd1 a_21740_17623# a_21652_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1760 vccd1 a_25660_7080# a_25572_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1761 a_22157_23336# a_14428_23544# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1762 vssd1 a_8454_21572# a_3703_18840# vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1763 a_5899_20244# a_5423_19668# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1764 a_14460_7080# a_14372_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1765 a_18380_9783# a_18292_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1766 a_1996_24328# a_7884_24328# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1767 a_13604_18884# a_5836_22760# vssd1 vssd1 nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1768 a_10296_13016# a_9744_13016# a_10092_13016# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1769 a_7804_9831# a_7496_9880# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1770 a_7259_24800# a_10452_18840# vssd1 vssd1 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1771 a_25212_8648# a_25124_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1772 a_20652_22424# a_20196_22112# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X1773 vssd1 a_11451_16488# a_5020_15796# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1774 vccd1 a_25648_25560# EOC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1775 a_25660_22327# a_25572_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1776 vccd1 a_27004_19624# a_26916_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1777 vccd1 a_12732_13440# a_12628_13484# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1778 vssd1 a_1692_18885# a_4628_23633# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
D58 a_1692_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1779 a_16588_8215# a_16500_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1780 vccd1 a_13077_22805# a_15940_22065# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1781 vccd1 a_5836_22760# a_4631_20408# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1782 a_6692_25560# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1783 a_8247_13397# a_8519_13836# a_8435_13397# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1784 a_15800_20540# a_13588_20535# a_14860_20807# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1785 vssd1 a_4815_20408# a_14736_20156# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1786 a_2588_5079# a_2500_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1787 vccd1 a_19500_20759# a_19412_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1788 vssd1 a_8456_23632# a_8352_23676# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1789 a_13188_21324# a_12020_21720# a_12984_21324# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1790 vssd1 a_10036_16532# a_10740_16532# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1791 a_11461_15748# a_11341_15704# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1792 vccd1 a_17484_14487# a_17396_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1793 a_7281_7142# a_1692_17302# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1794 vccd1 a_14796_9783# a_14708_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1795 a_11455_10348# a_10555_10216# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X1796 a_2876_19712# a_2568_19756# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1797 vssd1 a_4481_24757# a_12880_13884# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1798 a_19724_6647# a_19636_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1799 SDAC[6] a_1772_23544# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1800 a_27452_22760# a_27364_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1801 vssd1 a_7672_20453# a_1692_16488# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1802 a_11856_12700# a_9332_12695# a_11544_12700# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1803 a_25324_12919# a_25236_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1804 a_27116_5079# a_27028_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1805 vccd1 a_14796_6647# a_14708_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1806 a_3415_18885# a_1804_21723# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1807 a_19868_23588# a_9900_24756# a_19556_23992# vssd1 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1808 SDAC[5] a_1772_20408# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1809 a_8548_18884# a_4815_20408# a_11788_18884# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1810 vssd1 a_4573_17272# a_4693_17316# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1811 vssd1 a_11011_15704# a_10396_16488# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1812 a_21852_5512# a_21764_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1813 vccd1 a_27564_16055# a_27476_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1814 a_23196_8648# a_23108_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D59 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1815 vccd1 a_9420_6647# a_9332_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1816 vccd1 a_9900_24756# a_13508_23588# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1817 vccd1 a_16364_16055# a_16276_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1818 vccd1 a_27564_12919# a_27476_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1819 vccd1 a_1772_25112# SC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1820 vccd1 a_4481_24757# a_5627_23544# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X1821 a_12424_13484# a_11872_13467# a_12220_13484# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1822 vccd1 a_19276_5079# a_19188_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1823 a_4576_17020# a_2464_16603# a_4264_17020# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1824 vccd1 a_27564_8215# a_27476_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1825 vccd1 a_15804_11784# a_15716_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1826 a_21404_13352# a_21316_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1827 vccd1 a_19500_11351# a_19412_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1828 a_14544_21724# a_12020_21720# a_14232_21724# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1829 a_6643_15704# a_6973_15704# a_7093_16302# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1830 vssd1 a_10192_8692# a_4481_24757# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1831 a_21404_10216# a_21316_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1832 vssd1 a_4236_26254# a_2444_26249# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1833 vssd1 a_22771_24765# a_20776_24766# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1834 DIGITAL_OUT[3] a_18256_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1835 a_1692_3944# a_1604_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1836 vccd1 a_7281_7142# a_9180_14609# vccd1 pfet_06v0 ad=0.5913p pd=3.27u as=0.2847p ps=1.615u w=1.095u l=0.5u
X1837 a_12351_16620# a_11451_16488# vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1838 vccd1 a_5940_6390# a_6172_9432# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1839 vssd1 a_22157_23336# a_22277_23380# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1840 vccd1 a_23532_20759# a_23444_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1841 a_20732_3511# a_20644_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1842 a_14756_20856# a_13588_20535# a_14552_20856# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1843 a_4220_8736# a_3912_8780# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1844 a_5132_7564# a_5831_11000# a_5767_11045# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1845 vssd1 a_20652_22424# a_25648_25560# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1846 vccd1 a_1772_15704# SDAC[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1847 a_11548_13824# a_13496_15774# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1848 a_21392_25940# a_20196_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1849 a_14460_3511# a_14372_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1850 vccd1 a_1772_12568# SDAC[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1851 vccd1 a_13564_5512# a_13476_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1852 a_18268_5512# a_18180_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1853 vssd1 a_1692_26427# a_1604_26471# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1854 a_27900_21192# a_27812_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1855 a_14649_21584# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X1856 vccd1 a_20396_16055# a_20308_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1857 a_13653_24948# a_13533_24904# a_12909_24837# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1858 a_26108_19624# a_26020_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1859 a_17820_13352# a_17732_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1860 vccd1 a_24092_13352# a_24004_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1861 a_6006_18884# a_5530_18884# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1862 a_9211_17272# a_9559_17540# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X1863 vccd1 a_11011_15704# a_10396_16488# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1864 a_15371_24947# a_14895_24372# a_15119_24394# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1865 vssd1 a_1804_21723# a_1716_21767# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1866 a_8736_19363# a_1916_17302# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1867 vccd1 a_23532_14487# a_23444_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1868 a_21404_7080# a_21316_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1869 a_25324_9783# a_25236_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1870 a_5844_9880# a_5724_9432# vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X1871 a_17820_10216# a_17732_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1872 a_11760_11828# a_10787_11829# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1873 vccd1 a_27452_19624# a_27364_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1874 vccd1 a_1812_17353# a_5412_15495# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1875 vssd1 a_6547_11045# a_6543_12612# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1876 vccd1 a_23532_11351# a_23444_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1877 a_16576_23676# a_16428_23943# a_16408_23676# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1878 a_2564_18884# a_2444_18840# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
D60 vssd1 a_1692_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1879 a_11676_20452# a_9920_20096# a_9560_20452# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1880 vssd1 a_14089_13744# a_13984_13884# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1881 a_3816_18588# a_1604_18584# a_2876_18144# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1882 vssd1 a_1772_15704# SDAC[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1883 vccd1 a_9980_5512# a_9892_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1884 a_27900_11784# a_27812_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1885 a_14348_20856# a_14248_20686# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1886 a_9360_11132# a_7639_11459# a_8232_11390# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1887 vccd1 a_23532_5079# a_23444_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1888 a_16700_11784# a_16612_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1889 vccd1 a_9920_20096# a_8940_21590# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1890 a_3619_14136# a_3949_14136# a_4069_14180# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1891 a_11856_12700# a_9744_13016# a_11544_12700# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1892 a_25772_12919# a_25684_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1893 a_1772_23544# a_3564_23544# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1894 a_3619_11000# a_3949_11000# a_4069_11044# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1895 vccd1 a_12108_21664# a_12020_21720# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1896 a_1772_20408# a_3564_20408# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1897 vccd1 a_20620_18056# a_20532_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1898 vccd1 a_13004_8648# a_12916_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1899 vccd1 a_6172_5512# a_6084_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1900 vssd1 a_5612_23118# a_1916_22021# vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1901 vccd1 a_24640_25940# DIGITAL_OUT[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1902 a_20672_24860# a_18951_24416# a_19544_24416# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1903 a_12351_16620# a_11451_16488# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X1904 vssd1 a_8764_15749# a_10228_15793# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1905 a_20732_21192# a_20644_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1906 a_8736_19363# a_5836_22760# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1907 a_6440_18056# a_8156_17584# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1908 vccd1 a_1772_25112# SC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1909 vccd1 a_26108_22760# a_26020_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1910 a_27452_3944# a_27364_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1911 a_15692_6647# a_15604_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1912 vccd1 a_14796_8648# a_14708_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1913 vssd1 a_7628_20155# a_7540_20199# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1914 a_21852_13352# a_21764_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1915 a_23084_5079# a_22996_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1916 vccd1 a_5237_13397# a_5642_14180# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1917 a_16155_13880# a_10871_12268# a_13900_12568# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1918 a_15849_22804# a_15119_22826# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X1919 a_10866_20152# a_5836_22760# a_10662_20152# vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1920 vssd1 a_5972_17720# a_8841_15448# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1921 a_10808_13880# a_8721_14920# a_10808_13396# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1922 a_21852_10216# a_21764_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1923 a_18853_23379# a_18733_23269# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1924 vccd1 a_6499_21264# a_5895_21372# vccd1 pfet_06v0 ad=0.3975p pd=2.185u as=0.1521p ps=1.105u w=0.585u l=0.5u
X1925 a_6118_14180# a_5642_14180# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1926 a_10808_17662# a_10215_17731# a_11544_17404# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1927 a_5237_13397# a_4233_13744# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1928 a_16252_5512# a_16164_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1929 a_6508_5079# a_6420_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1930 a_4233_10608# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1931 a_6981_14986# a_6861_15429# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1932 a_3072_10564# a_9744_8392# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1933 vssd1 a_8752_8648# a_7404_9006# vssd1 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X1934 vccd1 a_23980_20759# a_23892_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1935 a_13416_19756# a_13015_19712# a_12359_19624# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
D61 a_1692_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1936 vccd1 a_26108_16488# a_26020_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1937 a_10296_13016# a_9332_12695# a_10092_13016# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1938 a_4481_24757# a_10192_8692# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1939 a_7032_24047# a_6631_24003# a_5975_23812# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1940 a_14895_22804# a_14271_22804# a_14727_22804# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1941 vccd1 a_1772_15704# SDAC[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1942 a_11548_13824# a_13496_15774# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1943 a_9560_20452# a_9920_20096# a_12104_20452# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1944 a_19804_24460# a_19352_24460# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X1945 vccd1 a_1772_12568# SDAC[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1946 vccd1 a_18716_3511# a_18628_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1947 a_6796_25511# a_6488_25560# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1948 a_5879_19668# a_5423_19668# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1949 vccd1 a_22300_19624# a_22212_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1950 a_8736_19363# a_1916_17302# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1951 a_9612_15704# a_8736_19363# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1952 a_14652_12605# a_14089_13744# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1953 a_6175_11045# a_3703_18840# a_5132_7564# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
D62 vssd1 a_2140_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1954 vccd1 a_19164_3944# a_19076_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1955 vccd1 a_20508_8648# a_20420_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1956 a_26556_19624# a_26468_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1957 vccd1 a_19948_17623# a_19860_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1958 a_16120_23992# a_15568_23992# a_15916_23992# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1959 vccd1 a_20508_5512# a_20420_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1960 vccd1 a_23980_14487# a_23892_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1961 vccd1 a_8076_6647# a_7988_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1962 a_20859_26424# a_7884_24328# a_1996_24328# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1963 a_15456_19368# a_14708_18100# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
D63 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1964 DIGITAL_OUT[2] a_17024_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1965 a_2564_18884# a_2892_18840# a_2544_19306# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1966 vccd1 a_23980_11351# a_23892_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1967 a_7717_16324# a_7597_15704# a_6973_15704# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1968 vssd1 a_1772_15704# SDAC[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1969 a_11961_12656# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1970 a_20620_12919# a_20532_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1971 a_19612_7080# a_19524_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1972 a_6299_7608# a_5831_11000# a_1772_11000# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1973 SDAC[6] a_1772_23544# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1974 a_15244_8215# a_15156_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1975 vccd1 a_19164_10216# a_19076_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1976 a_25660_8648# a_25572_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1977 a_5084_25560# a_4628_25248# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X1978 a_9732_21236# a_7259_24800# a_7628_20155# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1979 a_2904_11916# a_1940_12312# a_2700_11916# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1980 a_9744_8392# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1981 a_21292_9783# a_21204_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1982 vccd1 a_13452_9783# a_13364_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1983 a_17947_24328# a_18295_24328# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X1984 vccd1 a_27004_7080# a_26916_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1985 vccd1 a_13452_6647# a_13364_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1986 a_10111_17775# a_9211_17272# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X1987 vccd1 a_20508_13352# a_20420_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1988 vccd1 a_14576_25200# a_14471_25571# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1989 a_4094_22596# a_3954_21976# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X1990 vssd1 a_1772_6296# SDAC[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1991 a_7022_18884# a_6358_19378# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1992 a_4693_17892# a_4573_17272# a_3949_17272# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1993 vccd1 a_13496_17337# a_11628_18056# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1994 a_18716_16488# a_18628_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D64 vssd1 a_2444_24328# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1995 vccd1 a_24640_25940# DIGITAL_OUT[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1996 a_7093_15748# a_6973_15704# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1997 a_9532_19624# a_1916_17302# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1998 vssd1 a_1772_3160# SDAC[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1999 a_12395_15540# a_11919_14964# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2000 a_4693_14756# a_4573_14136# a_3949_14136# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2001 vccd1 a_1692_8215# a_1604_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D65 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2002 DIGITAL_OUT[1] a_13216_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2003 vccd1 a_26556_22760# a_26468_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2004 vssd1 a_7820_7564# a_7192_9710# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2005 DIGITAL_OUT[3] a_18256_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2006 a_22244_22424# a_21684_22020# a_22116_22020# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X2007 vccd1 a_7820_7564# a_7192_9710# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2008 vssd1 a_6643_15704# a_3887_18840# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2009 a_27564_5079# a_27476_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2010 a_21964_25560# a_21864_25390# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2011 vccd1 a_26220_8215# a_26132_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2012 a_9744_25560# a_9332_25239# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2013 vccd1 a_11628_18056# a_9800_18056# vccd1 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2014 a_10428_3944# a_10340_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2015 a_22636_6647# a_22548_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2016 vssd1 a_3999_21676# a_3935_21720# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2017 DIGITAL_OUT[0] a_9408_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2018 a_11544_25244# a_9332_25239# a_10604_25511# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2019 a_16428_23943# a_16120_23992# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2020 a_6154_19460# a_5530_18884# a_6006_18884# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2021 a_28012_12919# a_27924_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2022 vccd1 a_23196_10216# a_23108_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2023 a_4731_20872# a_4631_20408# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2024 vccd1 a_8456_23632# a_8352_23676# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2025 a_12073_23152# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2026 vccd1 a_26556_16488# a_26468_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2027 vccd1 a_2444_26249# COMP_CLK vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2028 vssd1 a_18403_18493# a_16773_18528# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2029 a_9408_25940# a_2052_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2030 a_21404_19624# a_21316_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2031 vccd1 a_19052_16055# a_18964_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2032 vccd1 a_1916_17302# a_10555_21267# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2033 a_9532_19624# a_9900_13396# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2034 vssd1 a_8519_13836# a_8721_14920# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2035 vccd1 a_22188_5079# a_22100_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2036 vssd1 a_2968_17317# a_2668_9132# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2037 vccd1 a_12220_5512# a_12132_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2038 a_14367_25615# a_13467_25112# vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2039 vccd1 a_12413_11000# a_12533_11620# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
D66 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2040 a_22748_16488# a_22660_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2041 vccd1 a_25212_10216# a_25124_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2042 a_9560_20452# a_7259_24800# a_2444_24328# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2043 vssd1 a_6719_16532# a_7195_17107# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2044 vssd1 a_5940_6390# a_6971_9176# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2045 a_2892_18840# a_10555_21267# a_12132_19288# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2046 vccd1 a_18716_8648# a_18628_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2047 vssd1 a_13252_22804# a_9900_24756# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2048 vssd1 a_4752_15704# a_2140_17302# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2049 a_13672_13884# a_11460_13880# a_12732_13440# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2050 a_19612_3511# a_19524_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2051 vccd1 a_21203_23197# a_19308_23544# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2052 vccd1 a_18716_5512# a_18628_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2053 a_10752_25244# a_10604_25511# a_10584_25244# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2054 vccd1 a_26220_23895# a_26132_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D67 vssd1 a_1692_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2055 a_3036_3944# a_2948_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2056 vccd1 a_26108_3944# a_26020_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2057 a_22476_25511# a_22168_25560# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2058 a_5636_9476# a_1996_11000# a_4965_14136# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2059 a_1772_23544# a_3564_23544# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2060 vccd1 a_26220_20759# a_26132_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2061 vccd1 a_6440_18056# a_1692_18528# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
D68 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2062 a_19724_8215# a_19636_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2063 vccd1 a_12152_10304# a_11960_10348# vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2064 vssd1 a_14895_22804# a_15371_23379# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2065 a_17368_23676# a_15156_23671# a_16428_23943# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2066 vssd1 a_12262_23544# a_5940_6390# vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2067 vccd1 a_16588_10216# a_16500_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2068 vccd1 a_6643_15704# a_3887_18840# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2069 a_13488_11000# a_8927_13836# vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X2070 vccd1 a_9800_18056# a_8156_17584# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2071 a_25772_9783# a_25684_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2072 a_22636_17623# a_22548_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2073 a_6266_14756# a_5642_14180# a_6118_14180# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2074 vccd1 a_4828_3944# a_4740_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2075 a_21852_7080# a_21764_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2076 vccd1 a_25100_25463# a_25012_25560# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2077 vssd1 a_1692_10688# a_1604_13880# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2078 vccd1 a_8076_5512# a_7988_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2079 vccd1 a_17932_9783# a_17844_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2080 DIGITAL_OUT[0] a_9408_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2081 vccd1 a_17932_6647# a_17844_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2082 vssd1 a_1772_25112# SC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2083 vccd1 a_11548_13824# a_13588_20535# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2084 vccd1 a_20956_13352# a_20868_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2085 vssd1 a_1692_10688# a_1604_10744# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2086 vccd1 a_23084_16055# a_22996_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2087 a_23868_3511# a_23780_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2088 a_17372_11784# a_17284_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2089 vccd1 a_13496_17337# a_11628_18056# vccd1 pfet_06v0 ad=0.428p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2090 a_7820_7564# a_8121_13016# a_9687_10744# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2091 vccd1 a_26220_14487# a_26132_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2092 vccd1 a_23084_12919# a_22996_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2093 a_20620_6647# a_20532_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2094 a_10787_11829# a_10871_12268# a_10807_12312# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2095 a_6859_26515# a_6383_25940# a_6607_25962# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2096 a_1692_18528# a_6440_18056# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X2097 a_15120_14584# a_8721_14920# vccd1 vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2098 vccd1 a_7167_13188# a_7623_13166# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2099 vccd1 a_23980_5079# a_23892_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2100 vccd1 a_26220_11351# a_26132_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2101 vccd1 a_1692_10688# a_2948_9176# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2102 a_13832_15424# a_14092_14920# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2103 vccd1 a_15020_11351# a_14932_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2104 a_14908_3944# a_14820_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2105 vccd1 a_13452_8648# a_13364_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2106 vccd1 a_21404_16488# a_21316_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2107 a_1772_6296# a_3564_6296# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2108 a_1772_3160# a_3564_3160# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2109 a_8153_25200# a_7736_25244# a_8529_25244# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2110 vccd1 a_20172_5079# a_20084_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2111 vccd1 a_27900_3944# a_27812_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2112 DIGITAL_OUT[2] a_17024_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2113 vccd1 a_12073_23152# a_11968_23292# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2114 vccd1 a_4752_15704# a_2140_17302# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2115 vccd1 a_1692_7080# a_1604_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2116 vssd1 a_6736_23632# a_6631_24003# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2117 a_18268_7080# a_18180_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2118 vccd1 a_4236_26254# a_2444_26249# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2119 a_9408_25940# a_2052_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2120 a_21852_19624# a_21764_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2121 vssd1 a_1772_12568# SDAC[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2122 a_4481_24757# a_10192_8692# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X2123 a_23420_21192# a_23332_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2124 a_11628_18056# a_13496_17337# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2125 vccd1 a_26668_5079# a_26580_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2126 a_7709_7864# a_4348_7909# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2127 vssd1 a_9295_22596# a_9771_22020# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2128 vccd1 a_16700_5512# a_16612_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2129 vccd1 a_9744_8392# a_3072_10564# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2130 a_15816_23822# a_15119_24394# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2131 a_24540_13352# a_24452_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2132 a_6956_5079# a_6868_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2133 a_24092_3944# a_24004_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2134 a_12856_16620# a_12560_16976# a_11799_16488# vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2135 a_1692_17302# a_10900_14964# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X2136 a_17036_6647# a_16948_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2137 vccd1 a_25660_10216# a_25572_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2138 a_24540_10216# a_24452_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2139 vccd1 a_10192_8692# a_4481_24757# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2140 a_18161_23676# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2141 a_3542_22242# a_3954_21976# a_4094_22596# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2142 vccd1 a_17820_16488# a_17732_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2143 a_13280_10748# a_11559_10304# a_12152_10304# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2144 a_8852_15704# a_9900_13396# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2145 a_26108_18056# a_26020_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2146 a_11376_17404# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2147 a_6643_15704# a_6973_15704# a_7093_15748# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2148 a_7516_3944# a_7428_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2149 vccd1 a_13467_25112# a_10732_24328# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2150 vccd1 a_6328_17342# a_1692_10688# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2151 a_21740_20759# a_21652_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2152 a_26108_14920# a_26020_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2153 vssd1 a_10472_14181# a_5724_9432# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2154 a_20672_24860# a_19056_24816# a_19544_24416# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
D69 a_5940_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2155 vccd1 a_20956_8648# a_20868_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2156 vccd1 a_27900_18056# a_27812_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2157 vssd1 a_17024_25940# DIGITAL_OUT[2] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2158 vccd1 a_20956_5512# a_20868_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2159 vccd1 a_21628_3511# a_21540_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2160 a_11685_14180# a_11565_14136# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2161 a_18828_12919# a_18740_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D70 a_2444_24328# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2162 a_21292_12919# a_21204_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2163 a_19556_23992# a_9900_24756# a_19408_23992# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X2164 vccd1 a_15356_3511# a_15268_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2165 a_11909_10030# a_11789_9432# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2166 DIGITAL_OUT[0] a_9408_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2167 vssd1 a_1772_25112# SC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2168 vssd1 a_11235_14136# a_9992_12846# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
D71 a_1804_21723# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2169 a_15692_8215# a_15604_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2170 vccd1 a_4481_24757# a_9744_8392# vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2171 a_21740_14487# a_21652_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2172 a_1692_5079# a_1604_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2173 a_8736_19363# a_10452_18840# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X2174 a_21740_11351# a_21652_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2175 a_12560_16976# a_11548_13824# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2176 a_2772_22892# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2177 a_11636_21236# a_5019_20408# a_11392_21236# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X2178 vssd1 a_10452_18840# a_7259_24800# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2179 vccd1 a_27452_7080# a_27364_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2180 a_4233_15312# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2181 vccd1 a_4828_5079# a_4740_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2182 a_26220_5079# a_26132_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2183 a_16252_7080# a_16164_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2184 a_9161_9520# a_8744_9564# a_9537_9564# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2185 vssd1 a_18312_22021# a_12636_21976# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2186 vccd1 a_21852_16488# a_21764_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2187 a_2016_10331# a_1604_10744# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2188 a_11215_12312# a_8940_21590# a_10787_11829# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2189 a_6271_22596# a_5647_22020# a_6103_22596# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2190 a_14708_18100# a_13776_18100# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2191 a_4609_15452# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2192 vssd1 a_4771_21192# a_4403_21582# vssd1 nfet_06v0 ad=0.14985p pd=1.145u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2193 a_27004_8648# a_26916_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2194 a_7984_24372# a_7884_24328# vccd1 vccd1 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2195 a_13416_19756# a_13120_20112# a_12359_19624# vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2196 a_18268_3511# a_18180_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2197 vccd1 a_10452_18840# a_7259_24800# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2198 a_15371_17016# a_8144_19288# a_2444_18840# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2199 vssd1 a_18256_25560# DIGITAL_OUT[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2200 vccd1 a_11076_24372# a_14271_22804# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2201 vccd1 a_5600_18101# a_8583_20856# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2202 vccd1 a_18380_5079# a_18292_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2203 a_23644_23291# a_23833_25200# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2204 a_10876_3944# a_10788_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2205 a_2772_13484# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2206 vccd1 a_17024_25940# DIGITAL_OUT[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2207 SDAC[5] a_1772_20408# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2208 a_10616_17775# a_10320_17360# a_9559_17540# vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2209 a_8744_9564# a_6532_9559# a_7804_9831# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2210 a_5137_24860# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2211 vccd1 a_3036_8215# a_2948_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2212 a_2772_10348# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2213 a_23833_25200# a_23416_25244# a_24209_25244# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2214 vccd1 a_16588_9783# a_16500_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2215 vccd1 a_26668_17623# a_26580_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2216 vccd1 a_16588_6647# a_16500_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2217 vssd1 a_13496_17337# a_11628_18056# vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2218 vccd1 a_19164_14920# a_19076_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2219 vccd1 a_5940_6390# a_1772_11000# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2220 DIGITAL_OUT[5] a_24640_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2221 vccd1 a_14895_22804# a_15351_22826# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2222 a_7531_12403# a_7055_11828# a_7279_11850# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2223 a_23644_5512# a_23556_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2224 vccd1 a_19164_11784# a_19076_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2225 vssd1 a_13216_25940# DIGITAL_OUT[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2226 a_19056_24816# a_12108_21664# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2227 a_26556_18056# a_26468_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2228 vssd1 a_6499_21264# a_6495_21724# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2229 a_11392_21236# a_11292_21192# vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2230 a_17372_5512# a_17284_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2231 a_19357_21768# a_17221_20453# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2232 vssd1 a_17452_20108# a_12860_21976# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2233 a_26556_14920# a_26468_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2234 a_4681_16880# a_4264_17020# a_5057_17020# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2235 vccd1 a_20060_3944# a_19972_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2236 a_17844_25560# a_17396_25201# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2237 vccd1 a_19612_13352# a_19524_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2238 vssd1 a_3564_12568# a_1772_12568# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2239 a_10180_11828# a_1692_17302# a_9920_11828# vccd1 pfet_06v0 ad=0.1736p pd=1.18u as=0.224p ps=1.36u w=0.56u l=0.5u
X2240 a_13120_20112# a_12108_21664# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2241 a_14176_17020# a_12455_16576# a_13048_16576# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2242 a_3212_11872# a_2904_11916# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2243 vccd1 a_14068_23992# a_14403_24328# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X2244 vccd1 a_7452_21280# a_7348_21324# vccd1 pfet_06v0 ad=0.22725p pd=1.91u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2245 vssd1 a_2588_21976# a_2500_22020# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2246 vssd1 a_3887_18840# a_3823_18885# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2247 a_3484_3944# a_3396_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2248 vccd1 a_26556_3944# a_26468_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2249 a_22524_3511# a_22436_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2250 vccd1 a_7988_19668# a_11348_22065# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2251 vssd1 a_5836_22760# a_14372_18884# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X2252 a_8048_25244# a_5524_25239# a_7736_25244# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
D72 vssd1 a_6388_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2253 vccd1 a_1692_18528# a_5524_25239# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2254 a_7154_14756# a_6470_14674# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X2255 vccd1 a_15356_5512# a_15268_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2256 a_16252_3511# a_16164_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2257 a_22636_8215# a_22548_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2258 vccd1 a_23196_14920# a_23108_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2259 a_21392_25940# a_20196_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2260 a_3404_24812# a_5836_22760# a_5732_22804# vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2261 vccd1 a_2588_21976# a_2500_22020# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2262 a_16217_20496# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2263 vccd1 a_3816_23292# a_4233_23152# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2264 vssd1 a_1692_18528# a_1604_20152# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
D73 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2265 a_9940_15448# a_1916_17302# a_9736_15448# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.1722p ps=1.24u w=0.82u l=0.6u
X2266 vccd1 a_23196_11784# a_23108_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2267 a_14708_18100# a_13776_18100# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2268 vccd1 a_10428_7080# a_10340_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2269 vccd1 a_22524_21192# a_22436_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2270 a_11664_10704# a_11548_13824# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2271 vccd1 a_7628_20155# a_7540_20199# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2272 a_25324_17623# a_25236_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2273 vssd1 a_9744_8392# a_3072_10564# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2274 a_27116_9783# a_27028_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2275 vccd1 a_17785_23632# a_17680_23676# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2276 a_16112_20540# a_13588_20535# a_15800_20540# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2277 a_13029_24394# a_12909_24837# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2278 vccd1 a_23644_13352# a_23556_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2279 a_3228_17317# a_3479_18840# a_3415_18885# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2280 vccd1 a_25212_14920# a_25124_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2281 vccd1 a_25212_11784# a_25124_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2282 a_10988_5079# a_10900_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2283 vccd1 a_17024_25940# DIGITAL_OUT[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2284 vccd1 a_25324_5079# a_25236_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2285 a_19648_21976# a_6553_24373# vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X2286 a_5612_5079# a_5524_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2287 vccd1 a_3072_10564# a_8492_11448# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2288 a_21404_14920# a_21316_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2289 DIGITAL_OUT[5] a_24640_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2290 vccd1 a_11544_25244# a_11961_25200# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2291 a_12108_21664# a_15456_19368# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X2292 a_10192_8692# a_7988_3608# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
D74 vssd1 a_1692_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2293 vssd1 a_4481_24757# a_11939_17020# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X2294 a_18380_14487# a_18292_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2295 vssd1 a_13216_25940# DIGITAL_OUT[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2296 vssd1 CLK a_13496_17337# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2297 a_4481_24757# a_10192_8692# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2298 a_1692_8648# a_1604_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2299 a_14736_20156# a_13120_20112# a_13608_19712# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2300 a_10676_16152# a_10228_15793# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2301 a_11544_12700# a_9744_13016# a_10604_12967# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2302 vccd1 a_17820_3511# a_17732_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2303 vssd1 a_5132_7564# a_3608_8736# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2304 a_23845_24372# a_23725_24904# a_23101_24837# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2305 a_3024_15452# a_2876_15008# a_2856_15452# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2306 vccd1 a_24540_3944# a_24452_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2307 a_17484_6647# a_17396_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2308 vccd1 a_5132_7564# a_3608_8736# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2309 vccd1 a_3036_7080# a_2948_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2310 a_7672_20453# a_7932_20453# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2311 vccd1 a_16588_8648# a_16500_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2312 a_24540_19624# a_24452_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2313 a_4576_17020# a_2052_17016# a_4264_17020# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2314 vssd1 a_21336_23589# a_4236_26254# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2315 a_11628_18056# a_13496_17337# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2316 a_27197_24904# a_23644_23291# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2317 a_19948_20759# a_19860_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2318 a_21653_22826# a_21533_23269# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2319 a_24092_11784# a_24004_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2320 a_7964_3944# a_7876_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2321 vccd1 a_14012_3511# a_13924_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2322 a_1792_16532# a_1692_16488# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2323 a_20620_8215# a_20532_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2324 vccd1 a_10732_24328# a_10576_24372# vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X2325 vccd1 a_22771_24765# a_20776_24766# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2326 a_13077_22805# a_12073_23152# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2327 a_14232_21724# a_12432_21307# a_13292_21280# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2328 a_17820_18056# a_17732_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2329 vccd1 a_17372_18056# a_17284_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2330 vccd1 a_23532_19191# a_23444_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2331 a_9612_15704# a_16773_18528# a_16709_18584# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2332 a_17820_14920# a_17732_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2333 a_12262_23544# a_2444_24328# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X2334 a_8972_15749# a_9123_17317# a_8764_15749# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.4137p ps=1.9u w=0.815u l=0.6u
X2335 a_21292_22327# a_21204_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2336 vccd1 a_20508_19191# a_20420_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2337 a_2444_26249# a_4236_26254# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2338 a_27116_23895# a_27028_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2339 a_11548_13824# a_13496_15774# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2340 a_27900_16488# a_27812_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2341 a_19948_11351# a_19860_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2342 vccd1 a_6563_11784# a_6431_11828# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2343 a_11628_18056# a_13496_17337# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2344 vccd1 a_14908_7080# a_14820_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2345 vccd1 a_11405_23544# a_11525_24164# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2346 a_22948_22020# a_22244_22424# vccd1 vccd1 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2347 vccd1 a_22972_21192# a_22884_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2348 vccd1 a_4752_7864# a_3564_15704# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2349 a_24640_25940# a_24004_22804# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2350 vccd1 a_12108_21664# a_21204_25239# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2351 a_23728_25244# a_21204_25239# a_23416_25244# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2352 a_25772_17623# a_25684_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2353 vccd1 a_5084_25560# a_13216_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D75 vssd1 a_1692_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2354 vccd1 a_20196_25940# a_21392_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2355 vssd1 a_3072_10564# a_10864_23292# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2356 vccd1 a_2444_24328# a_13252_22804# vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2357 a_5020_12613# a_8721_14920# vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X2358 a_7316_9176# a_1996_11000# a_6563_11784# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2359 vccd1 a_3564_9432# a_1772_9432# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2360 vccd1 a_25660_14920# a_25572_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2361 a_13280_10748# a_11664_10704# a_12152_10304# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2362 a_22476_25511# a_22168_25560# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2363 a_16744_22042# a_16388_22424# vccd1 vccd1 pfet_06v0 ad=0.4488p pd=2.92u as=0.458p ps=2.02u w=1.02u l=0.5u
X2364 vccd1 a_25212_22327# a_25124_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2365 vccd1 a_3564_6296# a_1772_6296# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2366 vccd1 a_3564_3160# a_1772_3160# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2367 a_24988_3511# a_24900_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2368 a_17036_8215# a_16948_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2369 vccd1 a_25660_11784# a_25572_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2370 vssd1 a_11405_23544# a_11525_23588# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2371 a_7605_13972# a_7485_13928# a_6861_13861# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2372 a_8121_13016# a_7391_12612# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2373 a_3036_5079# a_2948_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2374 a_27452_8648# a_27364_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2375 a_2588_21976# a_2918_21976# a_3038_22020# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2376 a_14953_22424# a_14223_22020# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2377 a_20060_13352# a_19972_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2378 a_21740_6647# a_21652_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2379 a_23084_9783# a_22996_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2380 vccd1 a_18716_10216# a_18628_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2381 EOC a_25648_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2382 a_11656_23292# a_9444_23288# a_10716_22848# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2383 a_18403_18493# a_18733_18565# a_18853_18122# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2384 vccd1 a_14652_12605# a_14538_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X2385 vccd1 a_15244_9783# a_15156_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2386 a_20060_10216# a_19972_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2387 a_6488_25560# a_5524_25239# a_6284_25560# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2388 vccd1 a_24540_16488# a_24452_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2389 a_21852_14920# a_21764_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2390 a_6981_13971# a_6861_13861# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2391 vccd1 a_24092_7080# a_24004_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2392 vssd1 a_1692_26427# a_8671_22020# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2393 a_16155_15448# a_5831_12568# a_6172_9432# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2394 vccd1 a_15244_6647# a_15156_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2395 vssd1 a_9263_20408# a_9199_20453# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2396 vssd1 a_2444_24328# a_16155_13880# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2397 vssd1 a_6266_10260# a_6742_10836# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2398 a_22300_5512# a_22212_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2399 a_5831_11000# a_7526_10282# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2400 vccd1 a_21292_5079# a_21204_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2401 vccd1 a_8940_21590# a_9479_10261# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2402 a_27900_22327# a_27812_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2403 DIGITAL_OUT[1] a_13216_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2404 a_4573_17272# a_2544_19306# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2405 vccd1 a_28012_8215# a_27924_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2406 a_18256_25560# a_17844_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2407 a_23555_23544# a_23885_23544# a_24005_24142# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2408 a_2772_22892# a_1604_23288# a_2568_22892# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2409 a_21740_19191# a_21652_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2410 vssd1 a_10192_8692# a_4481_24757# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2411 a_6047_19668# a_5423_19668# a_5899_20244# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2412 a_21740_16055# a_21652_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2413 a_24428_6647# a_24340_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2414 vccd1 a_17820_8648# a_17732_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2415 a_13616_17020# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2416 vccd1 a_4481_24757# a_9744_8392# vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2417 vccd1 a_5880_12288# a_1692_18885# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2418 vccd1 a_23555_23544# a_21864_25390# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2419 a_12432_21307# a_12020_21720# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2420 vccd1 a_16588_12919# a_16500_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2421 vccd1 a_17820_5512# a_17732_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D76 a_2444_24328# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2422 vccd1 a_19724_14487# a_19636_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2423 a_2140_3944# a_2052_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2424 vccd1 a_25212_3944# a_25124_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2425 vssd1 a_6239_11000# a_6175_11045# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2426 vccd1 a_22244_22424# a_22948_22020# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X2427 a_2052_19288# a_1604_18929# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2428 vccd1 a_23980_19191# a_23892_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2429 vccd1 a_22748_10216# a_22660_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2430 vccd1 a_5539_23589# a_5759_25940# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2431 a_6503_19690# a_6047_19668# a_6271_19690# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2432 a_2444_26249# a_4236_26254# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2433 a_27564_23895# a_27476_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2434 vccd1 a_4088_7909# a_3564_3160# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2435 vccd1 a_3932_3944# a_3844_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2436 a_1804_21723# a_12132_26424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X2437 vssd1 a_12073_23152# a_11968_23292# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X2438 a_12359_19624# a_13120_20112# a_12911_19756# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X2439 vccd1 a_18604_16055# a_18516_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2440 a_2772_13484# a_1604_13880# a_2568_13484# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2441 vccd1 a_14012_5512# a_13924_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2442 vccd1 a_7180_5512# a_7092_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2443 a_7820_7564# a_4964_9880# a_9479_10261# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2444 a_14455_22574# a_13999_22596# a_14223_22020# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2445 a_8568_7930# a_8752_8648# vccd1 vccd1 pfet_06v0 ad=0.4488p pd=2.92u as=0.458p ps=2.02u w=1.02u l=0.5u
X2446 a_11628_18056# a_13496_17337# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2447 a_2772_10348# a_1604_10744# a_2568_10348# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2448 a_22157_23336# a_14428_23544# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2449 a_22972_3511# a_22884_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2450 vccd1 a_1804_21723# a_4516_9521# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2451 a_2364_22892# a_2264_22848# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2452 a_11788_18884# a_10452_18840# a_8736_19363# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2453 a_10092_13016# a_9992_12846# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2454 a_20508_11784# a_20420_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2455 EOC a_25648_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2456 a_7259_24800# a_10452_18840# vccd1 vccd1 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2457 vssd1 a_13496_15774# a_11548_13824# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
D77 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2458 vccd1 a_20196_25940# a_21392_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2459 a_8791_20453# a_5940_6390# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2460 vssd1 a_17859_24373# a_19868_23588# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X2461 a_12108_21664# a_15456_19368# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2462 vssd1 a_12108_21664# a_21204_25239# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2463 vccd1 a_5500_13352# a_5412_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2464 vccd1 a_23196_3944# a_23108_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2465 vccd1 a_25660_22327# a_25572_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2466 vssd1 a_8156_17584# a_6328_17342# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2467 a_3220_16620# a_2052_17016# a_3016_16620# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2468 vssd1 a_9161_9520# a_9056_9564# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
D78 vssd1 a_5940_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2469 vccd1 a_10876_7080# a_10788_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2470 vccd1 a_22188_17623# a_22100_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2471 a_23644_7080# a_23556_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2472 a_27564_9783# a_27476_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2473 a_8009_11828# a_7279_11850# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2474 a_12911_19756# a_11787_20027# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.33755p ps=1.955u w=0.505u l=0.5u
X2475 a_7019_12612# a_6543_12612# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2476 vccd1 a_19724_9783# a_19636_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2477 vssd1 a_7055_11828# a_7531_12403# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2478 a_2544_19306# a_1996_11000# a_2564_18884# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2479 a_2364_13484# a_2264_13440# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2480 vccd1 a_19724_6647# a_19636_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2481 vccd1 a_25212_24328# a_25124_24372# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2482 a_11292_18884# a_4815_20408# a_8548_18884# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2483 SDAC[4] a_1772_15704# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2484 a_17372_7080# a_17284_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2485 a_7884_24328# a_9519_22020# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2486 a_11412_21720# a_4631_20408# a_11392_21236# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2487 a_2364_10348# a_2264_10304# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2488 vssd1 a_9900_24756# a_21684_22020# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2489 vccd1 a_25212_21192# a_25124_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2490 a_8736_19363# a_5836_22760# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X2491 a_10174_18884# a_5836_22760# a_9980_18884# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2492 a_28012_17623# a_27924_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2493 a_12720_10748# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2494 a_5767_11045# a_4964_9880# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2495 vccd1 a_23416_25244# a_23833_25200# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2496 vccd1 a_22636_16055# a_22548_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2497 vccd1 a_25772_5079# a_25684_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2498 a_9147_22020# a_8671_22020# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2499 vccd1 a_22636_12919# a_22548_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2500 vccd1 a_4569_12176# a_4464_12316# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2501 a_22168_25560# a_21204_25239# a_21964_25560# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2502 vccd1 a_9744_8392# a_3072_10564# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2503 a_16140_6647# a_16052_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2504 vccd1 a_7988_3608# a_10192_8692# vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2505 vssd1 a_4481_24757# a_13955_25236# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X2506 vccd1 a_15244_8648# a_15156_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2507 a_12262_23544# a_2444_24328# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X2508 vccd1 a_18403_21629# a_17452_20108# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2509 a_10616_20452# a_7259_24800# a_2444_24328# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2510 vccd1 a_10555_10216# a_8927_13836# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2511 a_14367_25615# a_13467_25112# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X2512 a_22412_23895# a_22324_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2513 vccd1 a_1692_18528# a_1604_23288# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2514 a_6620_3944# a_6532_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2515 vccd1 a_3484_7080# a_3396_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2516 SC a_1772_25112# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2517 vssd1 a_13533_24904# a_13653_24948# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2518 a_17024_25940# a_16388_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2519 vccd1 a_1916_22021# a_1828_22065# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2520 a_6098_14756# a_5642_14180# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2521 a_1692_10688# a_6328_17342# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2522 vccd1 a_20732_3511# a_20644_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2523 vssd1 a_4481_24757# a_16576_23676# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2524 vssd1 a_1692_10688# a_2948_9176# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2525 vccd1 a_14460_3511# a_14372_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2526 vssd1 a_3072_10564# a_7123_11124# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X2527 a_8748_5079# a_8660_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2528 a_4965_14136# a_5724_9432# a_5636_9476# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2529 vccd1 a_9900_24756# a_18996_23588# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2530 vccd1 a_1692_10688# a_1604_13880# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2531 a_10584_12700# a_9744_13016# a_10296_13016# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2532 a_20956_11784# a_20868_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2533 vssd1 a_1692_18528# a_1604_18584# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2534 SDAC[4] a_1772_15704# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2535 a_13832_15424# a_14092_14920# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2536 a_7535_11503# a_6635_11000# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X2537 EOC a_25648_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2538 a_4771_21192# a_5547_21551# a_5139_21292# vccd1 pfet_06v0 ad=0.1079p pd=0.935u as=0.1826p ps=1.71u w=0.415u l=0.5u
X2539 vssd1 a_1692_10688# a_1604_15448# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2540 SDAC[3] a_1772_12568# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2541 vccd1 a_13496_17337# a_11628_18056# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2542 a_17372_16488# a_17284_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2543 a_10599_11829# a_10871_12268# a_10787_11829# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2544 a_24629_24164# a_24509_23544# a_23885_23544# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2545 a_11292_21192# a_11324_19624# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2546 vccd1 a_26220_19191# a_26132_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2547 vccd1 a_3932_5079# a_3844_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2548 vccd1 a_3999_21676# a_5647_22020# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2549 vssd1 a_13494_14136# a_1916_17302# vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2550 vccd1 a_22748_8648# a_22660_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2551 DIGITAL_OUT[4] a_21392_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2552 a_19477_22804# a_19357_23336# a_18733_23269# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2553 vssd1 a_16217_20496# a_16112_20540# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X2554 a_2052_19288# a_1604_18929# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X2555 vccd1 a_2876_15008# a_2772_15052# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2556 vccd1 a_22748_5512# a_22660_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2557 a_17372_3511# a_17284_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2558 a_13272_21724# a_12432_21307# a_12984_21324# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2559 a_9744_25560# a_9332_25239# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2560 a_24629_23588# a_24509_23544# a_23885_23544# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2561 vccd1 a_25660_24328# a_25572_24372# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2562 a_18403_23197# a_18733_23269# a_18853_23379# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2563 a_22972_22760# a_22884_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2564 a_24540_24328# a_24452_24372# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2565 a_18268_13352# a_18180_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2566 a_17484_8215# a_17396_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2567 vccd1 a_25660_21192# a_25572_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2568 vccd1 a_5577_9040# a_5472_9180# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2569 a_18268_10216# a_18180_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2570 a_24005_23588# a_23885_23544# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2571 a_9956_21236# a_4815_20408# a_9732_21236# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2572 a_3484_5079# a_3396_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2573 a_3072_10564# a_9744_8392# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2574 vccd1 a_2140_8215# a_2052_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2575 a_14272_23992# a_13508_23588# a_14068_23992# vccd1 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2576 vccd1 a_2588_3944# a_2500_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2577 vccd1 a_15692_9783# a_15604_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2578 a_17844_25560# a_17396_25201# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X2579 vssd1 a_1692_18528# a_9444_23288# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2580 a_20060_19624# a_19972_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2581 vssd1 a_23555_23544# a_21864_25390# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2582 a_26668_20759# a_26580_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2583 a_28012_5079# a_27924_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2584 vccd1 a_15692_6647# a_15604_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2585 vccd1 a_6755_7864# a_6239_11000# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2586 a_13851_22020# a_13375_22020# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2587 a_3816_13884# a_2016_13467# a_2876_13440# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2588 vssd1 a_11324_19624# a_12132_26424# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2589 a_6047_19668# a_5423_19668# a_5879_19668# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2590 a_13019_15539# a_12543_14964# a_12767_14986# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2591 a_3816_10748# a_2016_10331# a_2876_10304# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2592 vccd1 a_19612_19191# a_19524_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2593 a_2568_15052# a_2016_15035# a_2364_15052# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2594 a_24092_8648# a_24004_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2595 a_22860_23895# a_22772_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2596 a_4731_20872# a_5019_20408# vccd1 vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2597 a_9744_13016# a_9332_12695# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2598 a_21516_18056# a_21428_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2599 vccd1 a_21068_18056# a_20980_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2600 a_24540_14920# a_24452_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2601 vssd1 a_4760_12613# a_4672_12657# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2602 vccd1 a_18256_25560# DIGITAL_OUT[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2603 a_22556_22020# a_9900_24756# a_22244_22424# vssd1 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2604 vssd1 a_12152_10304# a_11960_10348# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2605 a_19948_16055# a_19860_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2606 SDAC[3] a_1772_12568# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2607 a_1692_10688# a_6328_17342# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2608 a_12668_3944# a_12580_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2609 a_26668_14487# a_26580_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2610 vssd1 a_10192_8692# a_4481_24757# vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2611 a_9161_9520# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2612 a_12482_11828# a_12026_11828# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2613 a_24876_6647# a_24788_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2614 a_26668_11351# a_26580_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2615 vccd1 a_9920_20096# a_9444_19668# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2616 a_15468_11351# a_15380_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2617 a_11459_11000# a_11789_11000# a_11909_11598# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2618 vccd1 a_25660_3944# a_25572_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2619 a_7167_13188# a_6543_12612# a_7019_12612# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2620 a_17036_12919# a_16948_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2621 a_21292_17623# a_21204_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2622 a_7175_16554# a_6719_16532# a_6943_16554# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2623 a_2444_26249# a_4236_26254# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2624 vssd1 a_8492_24328# a_8444_24856# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X2625 a_7524_8692# a_7404_9006# vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X2626 a_4698_22596# a_4578_21976# a_3954_21976# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2627 a_4388_19288# a_1916_17302# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X2628 vccd1 a_18716_14920# a_18628_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2629 vccd1 a_19276_12919# a_19188_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2630 a_10555_21267# a_9900_13396# a_10759_21720# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X2631 vccd1 a_14460_5512# a_14372_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2632 a_19164_5512# a_19076_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2633 a_21740_8215# a_21652_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2634 vccd1 a_18716_11784# a_18628_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2635 vccd1 a_4771_21192# a_4403_21582# vccd1 pfet_06v0 ad=0.3276p pd=1.62u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2636 vccd1 a_4573_17272# a_4693_17892# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2637 a_12413_11000# a_8927_13836# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2638 vccd1 a_4573_14136# a_4693_14756# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2639 a_12543_14964# a_11919_14964# a_12395_15540# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2640 a_16140_10216# a_16052_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2641 a_8800_11132# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2642 vssd1 a_6553_24373# a_6431_22804# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2643 vccd1 a_1692_18528# a_9444_23288# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2644 a_4233_20016# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2645 a_2016_18171# a_1604_18584# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2646 vccd1 a_10396_16488# a_10240_16532# vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X2647 vssd1 a_9540_12268# a_4492_18840# vssd1 nfet_06v0 ad=0.224p pd=1.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2648 vccd1 a_9532_19624# a_9444_19668# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X2649 vccd1 a_20060_16488# a_19972_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2650 a_22300_7080# a_22212_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2651 a_26220_9783# a_26132_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2652 vccd1 a_1692_10688# a_6532_9559# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2653 a_5237_18101# a_4233_18448# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2654 a_2016_15035# a_1604_15448# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2655 a_5276_3944# a_5188_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D79 vssd1 a_1692_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2656 a_5769_24856# a_4481_24757# a_5137_24860# vssd1 nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
X2657 vssd1 a_11628_18056# a_9800_18056# vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2658 a_19544_24416# a_18951_24416# a_20280_24860# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2659 vssd1 a_3564_23544# a_1772_23544# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2660 vssd1 a_11279_12268# a_11215_12312# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2661 vccd1 a_3703_18840# a_3207_19288# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2662 a_6266_14756# a_5642_14180# a_6098_14756# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2663 a_7709_7864# a_4348_7909# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2664 a_2672_21782# a_2820_21192# a_2672_21237# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X2665 a_17632_21976# a_16388_22424# vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X2666 a_23420_22327# a_23332_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2667 a_14544_21724# a_12432_21307# a_14232_21724# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2668 a_24428_8215# a_24340_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2669 vccd1 a_9408_25940# DIGITAL_OUT[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2670 vssd1 a_5940_6390# a_15371_17016# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2671 a_12412_10348# a_11960_10348# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X2672 SC a_1772_25112# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2673 vccd1 a_7672_20453# a_1692_16488# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2674 a_2772_18188# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2675 vccd1 a_22748_14920# a_22660_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2676 a_10095_10744# a_8940_21590# a_7820_7564# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2677 a_24509_23544# a_22948_22020# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2678 vccd1 a_22636_9783# a_22548_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2679 vccd1 a_14708_18100# a_13496_15774# vccd1 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2680 a_1872_14602# a_1772_14136# vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2681 vccd1 a_22748_11784# a_22660_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2682 vssd1 a_6440_18056# a_1692_18528# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2683 vccd1 a_22636_6647# a_22548_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2684 vccd1 a_19164_19624# a_19076_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2685 a_21964_18056# a_21876_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2686 a_25212_22760# a_25124_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2687 vccd1 a_7988_3608# a_10192_8692# vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2688 a_8940_21590# a_9920_20096# a_11669_24856# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2689 vccd1 a_6266_14756# a_6702_14756# vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2690 vccd1 a_2140_7080# a_2052_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2691 vssd1 a_9800_18056# a_8156_17584# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2692 vccd1 a_2588_5079# a_2500_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2693 vccd1 a_15692_8648# a_15604_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2694 vssd1 a_1916_17302# a_8756_18884# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2695 a_4815_20408# a_9920_20096# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2696 vssd1 a_4481_24757# a_10752_25244# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
D80 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2697 a_24509_23544# a_22948_22020# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2698 vccd1 a_25324_16055# a_25236_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2699 a_19612_11784# a_19524_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2700 vccd1 a_25324_12919# a_25236_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2701 vccd1 a_27116_5079# a_27028_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2702 vccd1 a_8636_7080# a_8548_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D81 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2703 a_17484_12919# a_17396_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2704 a_7404_5079# a_7316_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2705 a_7744_11088# a_1692_10688# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2706 a_7597_15704# a_4716_18840# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2707 a_9687_10744# a_4964_9880# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2708 a_7001_19668# a_6271_19690# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2709 a_18847_24460# a_17947_24328# vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2710 a_9980_18884# a_1916_17302# vssd1 vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2711 a_17932_14487# a_17844_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2712 a_11961_12656# a_11544_12700# a_12337_12700# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2713 a_3072_10564# a_9744_8392# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X2714 a_10807_12312# a_7988_19668# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2715 a_19352_24460# a_19056_24816# a_18295_24328# vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2716 a_23555_23544# a_23885_23544# a_24005_23588# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2717 vssd1 a_5237_19669# a_5759_20452# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2718 vssd1 a_6047_19668# a_6523_20243# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2719 vccd1 a_19612_3511# a_19524_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2720 a_2364_13484# a_2264_13440# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2721 a_3220_16620# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2722 vssd1 a_10900_14964# a_1692_17302# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2723 a_19276_6647# a_19188_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2724 a_2364_10348# a_2264_10304# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2725 vssd1 a_6383_25940# a_6859_26515# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2726 vccd1 a_5795_21280# a_5547_21551# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2727 vccd1 a_21404_8648# a_21316_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2728 a_26108_5512# a_26020_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2729 vccd1 a_23196_19624# a_23108_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2730 vccd1 a_4815_20408# a_9076_15704# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2731 vssd1 a_8156_17584# a_6440_18056# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2732 vccd1 a_21404_5512# a_21316_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2733 vssd1 a_19056_24816# a_18951_24416# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2734 vccd1 a_8156_17584# a_6328_17342# vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2735 vssd1 a_12543_14964# a_13019_15539# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
D82 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
D83 vssd1 a_1804_21723# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2736 vccd1 a_1772_9432# SDAC[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2737 a_12888_10748# a_11960_10348# a_12720_10748# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2738 vssd1 a_20776_24766# a_20672_24860# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2739 vccd1 a_1772_6296# SDAC[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2740 a_23644_11784# a_23556_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2741 vccd1 a_27900_10216# a_27812_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2742 vccd1 a_1772_3160# SDAC[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2743 vccd1 a_23868_3511# a_23780_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2744 a_4828_5512# a_4740_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2745 a_16140_8215# a_16052_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2746 a_8972_15749# a_8852_15704# a_8764_15749# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2747 vccd1 a_20620_9783# a_20532_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2748 vssd1 a_17844_25560# a_18256_25560# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2749 a_2140_5079# a_2052_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2750 vccd1 a_20652_22424# a_25648_25560# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2751 vccd1 a_25212_19624# a_25124_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2752 a_7666_18884# a_7190_18884# a_7414_18884# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2753 a_9572_18884# a_5836_22760# a_8548_18884# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2754 vccd1 a_20620_6647# a_20532_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2755 a_11909_11044# a_11789_11000# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2756 vccd1 a_9408_25940# DIGITAL_OUT[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2757 vssd1 a_15392_13824# a_8519_13836# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
D84 vssd1 a_1692_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2758 vccd1 a_15064_25502# a_14872_25615# vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2759 a_4578_21976# a_4315_21237# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2760 a_7736_25244# a_5936_25560# a_6796_25511# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2761 vccd1 a_9800_18056# a_8156_17584# vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2762 vssd1 a_11459_11000# a_11279_12268# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
D85 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2763 a_8644_14181# a_6388_6390# a_8624_14602# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.4137p ps=1.9u w=0.815u l=0.6u
X2764 a_8736_25940# a_2500_22020# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2765 a_8752_8648# a_9161_9520# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2766 a_13496_17337# CLK vccd1 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2767 vssd1 a_4481_24757# a_6944_25244# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2768 a_25660_22760# a_25572_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2769 a_3642_22596# a_3542_22242# a_2918_21976# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2770 vccd1 a_13776_18100# a_14708_18100# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2771 a_13308_16620# a_12856_16620# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X2772 a_23532_12919# a_23444_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2773 a_3816_23292# a_2016_22875# a_2876_22848# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2774 a_4128_23292# a_2016_22875# a_3816_23292# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2775 vssd1 a_1772_20408# SDAC[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2776 vssd1 a_10555_10216# a_8927_13836# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2777 a_11544_17404# a_10616_17775# a_11376_17404# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2778 vccd1 a_25772_16055# a_25684_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2779 a_15800_20540# a_14000_20856# a_14860_20807# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2780 a_3816_20156# a_2016_19739# a_2876_19712# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2781 a_2352_11899# a_1940_12312# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2782 a_11324_3944# a_11236_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2783 a_27900_5512# a_27812_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2784 a_18853_21258# a_18733_21701# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2785 vccd1 a_25772_12919# a_25684_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2786 a_23532_6647# a_23444_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2787 a_8156_17584# a_9800_18056# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2788 vccd1 a_17036_9783# a_16948_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2789 vccd1 a_8232_11390# a_8040_11503# vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2790 a_9164_18884# a_1916_17302# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2791 DIGITAL_OUT[3] a_18256_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2792 a_14727_22804# a_14271_22804# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2793 a_11235_14136# a_11565_14136# a_11685_14180# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
D86 vssd1 a_5940_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2794 vccd1 a_17036_6647# a_16948_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2795 a_10576_24372# a_9812_24856# a_10372_24372# vccd1 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
D87 vssd1 XRST diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2796 vssd1 a_7988_3608# a_10192_8692# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2797 a_24092_16488# a_24004_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2798 vssd1 a_4752_7864# a_3564_15704# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2799 vccd1 a_2876_19712# a_2772_19756# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2800 DIGITAL_OUT[2] a_17024_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2801 a_24204_18056# a_24116_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2802 a_7778_14180# a_7302_14180# a_7526_14180# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2803 a_4128_13884# a_2016_13467# a_3816_13884# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
D88 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2804 vccd1 a_23084_5079# a_22996_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2805 a_8336_24372# a_7572_24856# a_8132_24372# vccd1 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
D89 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2806 a_4128_10748# a_2016_10331# a_3816_10748# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2807 a_9900_24756# a_13252_22804# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X2808 vccd1 a_21740_20759# a_21652_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2809 a_10604_12967# a_10296_13016# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2810 vccd1 a_7852_9006# a_6563_11784# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X2811 a_18156_11351# a_18068_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2812 a_5573_11829# a_4569_12176# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2813 vccd1 a_6508_5079# a_6420_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2814 vssd1 a_9744_8392# a_3072_10564# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2815 vccd1 a_19612_8648# a_19524_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2816 vccd1 a_19612_5512# a_19524_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2817 vccd1 a_18256_25560# DIGITAL_OUT[3] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2818 a_4264_17020# a_2464_16603# a_3324_16576# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2819 vccd1 a_27004_3944# a_26916_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2820 vssd1 a_22244_22424# a_22948_22020# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2821 vccd1 a_21180_21192# a_21092_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2822 vccd1 a_5612_23118# a_7706_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X2823 vccd1 a_18268_16488# a_18180_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2824 a_4760_12613# a_5020_12613# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2825 vssd1 a_21203_23197# a_19308_23544# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
D90 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2826 vssd1 a_13496_17337# a_11628_18056# vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2827 a_2568_19756# a_2016_19739# a_2364_19756# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2828 vccd1 a_21740_14487# a_21652_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2829 a_13999_22596# a_13375_22020# a_13851_22020# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2830 vccd1 a_25660_19624# a_25572_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2831 a_22188_20759# a_22100_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2832 vccd1 a_10740_16532# a_11936_17404# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2833 vccd1 a_21740_11351# a_21652_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2834 a_27004_13352# a_26916_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2835 vccd1 a_5724_3944# a_5636_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2836 a_6563_11784# a_7404_9006# a_7316_9176# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2837 a_27004_10216# a_26916_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2838 a_8764_15749# a_9076_15704# a_8972_15749# vssd1 nfet_06v0 ad=0.4137p pd=1.9u as=0.2119p ps=1.335u w=0.815u l=0.6u
D91 vssd1 a_2444_24328# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2839 a_26668_19191# a_26580_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2840 vccd1 a_2892_18840# a_2788_19288# vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2841 a_20060_14920# a_19972_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2842 a_13496_17337# CLK vccd1 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2843 a_26668_16055# a_26580_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2844 vccd1 a_20620_12919# a_20532_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2845 vssd1 a_4481_24757# a_9744_8392# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2846 vccd1 a_13900_8215# a_13812_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2847 a_6981_15539# a_6861_15429# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2848 a_23980_12919# a_23892_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2849 vccd1 a_18268_3511# a_18180_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2850 SDAC[6] a_1772_23544# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2851 a_24876_8215# a_24788_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2852 SDAC[5] a_1772_20408# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2853 vssd1 a_5940_6390# a_16155_15448# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2854 a_22188_14487# a_22100_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2855 vccd1 a_11324_19624# a_12132_26424# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X2856 vssd1 a_18984_22021# a_3564_23544# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2857 a_22188_11351# a_22100_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2858 a_10372_24372# a_9812_24856# a_10244_24856# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X2859 a_15804_3944# a_15716_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2860 vccd1 a_12668_7080# a_12580_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2861 a_11436_5079# a_11348_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2862 a_12413_11000# a_8927_13836# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2863 a_13216_25940# a_5084_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2864 vccd1 a_25648_25560# EOC vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2865 vccd1 a_24316_22760# a_24228_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2866 vccd1 a_9920_20096# a_2444_24328# vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2867 vssd1 a_4481_24757# a_22624_25244# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2868 a_8132_24372# a_7572_24856# a_8004_24856# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X2869 a_19164_7080# a_19076_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2870 DIGITAL_OUT[4] a_21392_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2871 vccd1 a_9532_13685# a_9444_13880# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X2872 vccd1 a_14649_21584# a_5836_22760# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2873 a_4041_24812# a_3728_24460# vccd1 vccd1 pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X2874 a_8144_19288# a_7414_18884# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2875 a_2140_8648# a_2052_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2876 vccd1 a_27564_5079# a_27476_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2877 a_2016_19739# a_1604_20152# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2878 vccd1 a_2968_17317# a_2668_9132# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2879 a_7852_5079# a_7764_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2880 a_6284_25560# a_2096_24372# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2881 a_5544_7584# a_5573_11829# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2882 vccd1 a_28012_16055# a_27924_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2883 a_7302_14180# a_6470_14674# a_7154_14756# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2884 vccd1 a_3703_18840# a_5559_13016# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2885 vccd1 a_28012_12919# a_27924_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2886 a_2772_18188# a_1604_18584# a_2568_18188# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2887 a_13496_17337# CLK vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2888 a_20060_5512# a_19972_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2889 a_2364_22892# a_2264_22848# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2890 a_8412_3944# a_8324_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2891 a_20508_16488# a_20420_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2892 a_2364_19756# a_1792_16532# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2893 vssd1 a_7337_25940# a_2820_21192# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2894 vccd1 a_4233_15312# a_4128_15452# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2895 a_14348_20856# a_14248_20686# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
D92 COMP_OUT vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2896 vssd1 a_13496_17337# a_11628_18056# vssd1 nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2897 vccd1 a_21852_8648# a_21764_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2898 vssd1 a_13048_16576# a_12856_16620# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2899 vccd1 a_21852_5512# a_21764_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2900 vccd1 a_22524_3511# a_22436_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2901 a_26556_5512# a_26468_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2902 a_17024_25940# a_16388_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2903 a_7452_21280# a_8736_25940# a_8791_20453# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2904 a_22188_6647# a_22100_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2905 a_27452_13352# a_27364_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2906 vccd1 a_16252_3511# a_16164_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2907 vssd1 a_12108_21664# a_12020_21720# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
D93 vssd1 a_2220_24686# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2908 vccd1 a_17372_10216# a_17284_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2909 a_27452_10216# a_27364_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D94 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2910 a_7623_13166# a_7167_13188# a_7391_12612# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2911 a_5975_23812# a_6736_23632# a_6527_24047# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X2912 a_5831_12568# a_7526_14180# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2913 a_2364_18188# a_2264_18144# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2914 a_3016_16620# a_2052_17016# a_2812_16620# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2915 vccd1 a_1692_3944# a_1604_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2916 a_3038_22574# a_2918_21976# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2917 vccd1 a_5836_22760# a_2444_24328# vccd1 pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2918 a_8736_19363# a_10452_18840# a_11292_18884# vssd1 nfet_06v0 ad=0.4161p pd=1.905u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2919 a_6887_11828# a_6431_11828# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2920 a_11787_20027# a_12359_19624# vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2921 vccd1 a_13496_17337# a_11628_18056# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2922 a_25436_3511# a_25348_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D95 a_2444_24328# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2923 vssd1 a_4088_7909# a_3564_3160# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2924 vccd1 a_24004_22804# a_24640_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2925 vccd1 a_23725_24904# a_23845_24372# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2926 vccd1 a_7337_25940# a_2820_21192# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2927 a_13216_25940# a_5084_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2928 vccd1 a_18268_8648# a_18180_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D96 vssd1 a_5940_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2929 a_19164_3511# a_19076_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2930 vssd1 a_15456_19368# a_12108_21664# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2931 a_3479_18840# a_6943_16554# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2932 vssd1 a_2140_17302# a_5020_12613# vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2933 vccd1 a_18268_5512# a_18180_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2934 vssd1 a_11760_11828# a_13280_10748# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2935 a_21203_23197# a_21533_23269# a_21653_22826# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2936 a_12780_21324# a_11392_21236# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2937 a_19276_8215# a_19188_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D97 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2938 a_11405_23544# a_2672_21782# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2939 a_16709_18584# a_8736_19363# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2940 vccd1 a_18380_14487# a_18292_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2941 a_11772_3944# a_11684_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2942 a_4964_9880# a_4516_9521# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2943 a_26220_12919# a_26132_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2944 a_23980_6647# a_23892_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2945 a_1772_23544# a_3564_23544# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2946 a_26108_7080# a_26020_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2947 vccd1 a_17484_9783# a_17396_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2948 a_10428_11351# a_10340_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2949 a_6776_25244# a_5936_25560# a_6488_25560# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2950 a_3004_21664# a_7259_24800# a_7175_24856# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X2951 a_13029_24947# a_12909_24837# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2952 vccd1 a_28012_24328# a_27924_24372# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2953 a_1772_20408# a_3564_20408# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2954 vssd1 a_13776_18100# a_14708_18100# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2955 a_15064_12613# a_14350_13016# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
D98 a_2140_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2956 vssd1 a_5612_17317# a_5524_17361# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2957 vccd1 a_17484_6647# a_17396_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2958 vccd1 a_27900_14920# a_27812_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2959 a_10555_10216# a_10903_10216# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X2960 a_11392_21236# a_5019_20408# a_11412_21720# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2961 vccd1 a_17260_16055# a_17172_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2962 vssd1 a_5020_15796# a_9532_13685# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2963 a_4752_7864# a_4716_18840# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X2964 a_15392_13824# a_14652_12605# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X2965 a_24540_5512# a_24452_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2966 vccd1 a_27900_11784# a_27812_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2967 vccd1 a_19948_20759# a_19860_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2968 a_2812_16620# a_2712_16576# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2969 vssd1 a_5539_23589# a_5759_25940# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2970 a_20172_6647# a_20084_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2971 vccd1 a_16700_11784# a_16612_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2972 a_22300_13352# a_22212_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2973 vccd1 a_26108_13352# a_26020_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2974 a_7952_9564# a_7804_9831# a_7784_9564# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2975 a_20956_16488# a_20868_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2976 a_5412_18101# a_1692_17302# a_5600_18101# vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2977 a_22300_10216# a_22212_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2978 vccd1 a_17844_25560# a_18256_25560# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2979 a_2444_24328# a_7259_24800# a_9560_20452# vssd1 nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2980 vssd1 a_10740_16532# a_11936_17404# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2981 vccd1 a_6956_5079# a_6868_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2982 a_26668_6647# a_26580_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2983 vssd1 a_9744_8392# a_3072_10564# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2984 vccd1 a_21292_22327# a_21204_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2985 a_10884_18884# a_10452_18840# a_8736_19363# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2986 vccd1 a_9800_14181# a_2220_11000# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2987 a_10871_12268# a_13910_11850# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2988 vccd1 a_19056_24816# a_18951_24416# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
D99 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2989 a_4380_3944# a_4292_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2990 vccd1 a_27452_3944# a_27364_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2991 vssd1 a_6755_7864# a_6239_11000# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2992 SDAC[6] a_1772_23544# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2993 vssd1 a_7485_13928# a_7605_13972# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2994 a_3912_8780# a_2948_9176# a_3708_8780# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2995 vssd1 a_8300_8648# a_8849_10744# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2996 a_11548_13824# a_13496_15774# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2997 vccd1 a_14796_10216# a_14708_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2998 vccd1 a_19948_11351# a_19860_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2999 vssd1 a_16388_25940# a_17024_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3000 a_9199_20453# a_5600_18101# a_7452_21280# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3001 vccd1 a_16428_23943# a_16324_23992# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3002 a_23420_3511# a_23332_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3003 a_13900_5079# a_13812_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3004 vssd1 a_4233_15312# a_4128_15452# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3005 a_27900_7080# a_27812_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3006 a_11459_9432# a_11789_9432# a_11909_9476# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
D100 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3007 COMP_CLK a_2444_26249# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3008 a_3935_21720# a_3703_18840# a_3507_21237# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3009 a_5076_23992# a_4628_23633# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3010 a_6103_22596# a_5647_22020# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3011 a_5159_21720# a_4403_21582# vssd1 vssd1 nfet_06v0 ad=48.6f pd=0.645u as=0.14985p ps=1.145u w=0.405u l=0.6u
X3012 a_18268_14920# a_18180_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3013 vccd1 a_16252_5512# a_16164_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3014 a_23532_8215# a_23444_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3015 vccd1 a_9744_8392# a_3072_10564# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3016 vssd1 a_7852_9006# a_7316_9176# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3017 a_27004_19624# a_26916_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3018 vccd1 a_21292_16055# a_21204_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3019 vccd1 a_18828_12919# a_18740_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3020 a_2016_22875# a_1604_23288# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
D101 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3021 vccd1 a_18312_22021# a_12636_21976# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3022 vccd1 a_21292_12919# a_21204_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3023 vccd1 a_24988_3511# a_24900_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3024 vccd1 a_11324_7080# a_11236_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3025 a_3304_17020# a_2464_16603# a_3016_16620# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3026 vccd1 a_21740_9783# a_21652_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3027 a_10092_25560# a_8836_24372# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3028 vssd1 a_25648_25560# EOC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3029 vccd1 a_15288_22021# a_14248_20686# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3030 a_9800_14181# a_8624_14602# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X3031 a_28012_9783# a_27924_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3032 vssd1 a_15456_19368# a_12108_21664# vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3033 a_3816_18588# a_2016_18171# a_2876_18144# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3034 vssd1 a_1772_15704# SDAC[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3035 vccd1 a_21740_6647# a_21652_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3036 a_7068_3944# a_6980_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3037 a_23725_24904# a_20260_23588# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3038 vccd1 a_1692_5079# a_1604_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D102 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3039 vssd1 a_10320_17360# a_10215_17731# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3040 a_13784_17020# a_12856_16620# a_13616_17020# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3041 a_11884_5079# a_11796_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3042 a_18156_16055# a_18068_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3043 a_14576_25200# a_12108_21664# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3044 vccd1 a_26220_5079# a_26132_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D103 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3045 a_10532_15448# a_1916_17302# a_10348_15448# vssd1 nfet_06v0 ad=0.1148p pd=1.1u as=0.1312p ps=1.14u w=0.82u l=0.6u
D104 vssd1 a_6388_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3046 vccd1 a_4220_8736# a_4116_8780# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3047 a_3527_21720# a_2164_21236# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3048 vccd1 a_27900_22327# a_27812_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3049 a_4128_13884# a_1604_13880# a_3816_13884# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
D105 a_1692_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3050 vccd1 a_24640_25940# DIGITAL_OUT[5] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3051 a_22116_22020# a_17859_24373# vssd1 vssd1 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3052 vccd1 a_13999_22596# a_14455_22574# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3053 a_10092_13016# a_9992_12846# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3054 vccd1 a_24428_9783# a_24340_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3055 a_4128_10748# a_1604_10744# a_3816_10748# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
D106 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3056 vccd1 a_1772_25112# SC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3057 a_2096_24372# a_1996_24328# vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3058 vccd1 a_27004_22760# a_26916_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3059 vccd1 a_24428_6647# a_24340_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3060 vccd1 a_26556_13352# a_26468_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3061 a_22456_25244# a_21616_25560# a_22168_25560# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
D107 vssd1 a_2220_24686# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3062 a_12449_23292# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3063 vccd1 a_24428_17623# a_24340_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3064 a_14392_14181# a_5972_17720# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X3065 a_2876_13440# a_2568_13484# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3066 vccd1 a_10451_23544# a_8456_23632# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3067 vssd1 a_17785_23632# a_17680_23676# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3068 a_18380_6647# a_18292_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3069 a_2876_10304# a_2568_10348# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3070 vssd1 a_9920_20096# a_13375_22020# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X3071 a_2444_24328# a_7259_24800# vccd1 vccd1 pfet_06v0 ad=0.52205p pd=2.045u as=0.4334p ps=2.85u w=0.985u l=0.5u
X3072 a_2588_21976# a_2918_21976# a_3038_22574# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3073 a_14428_23544# a_17785_23632# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3074 a_25212_5512# a_25124_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3075 a_13984_13884# a_11460_13880# a_13672_13884# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3076 vssd1 a_13120_20112# a_13015_19712# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3077 vccd1 a_27004_16488# a_26916_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3078 a_8860_3944# a_8772_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3079 a_13533_24904# a_4716_25204# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3080 a_9532_19624# a_9900_13396# a_9940_15448# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3081 a_7758_14734# a_7302_14180# a_7526_14180# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3082 a_22188_19191# a_22100_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3083 vccd1 a_1772_15704# SDAC[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3084 vssd1 a_16388_25940# a_17024_25940# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3085 a_17221_20453# a_16217_20496# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3086 vccd1 a_3072_10564# a_11068_17720# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3087 a_22188_16055# a_22100_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3088 vccd1 a_1772_12568# SDAC[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3089 vccd1 a_10428_3944# a_10340_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3090 a_7700_9880# a_6532_9559# a_7496_9880# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3091 vccd1 a_22972_3511# a_22884_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3092 a_3932_5512# a_3844_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3093 vccd1 a_12158_11784# a_12026_11828# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3094 a_10599_11829# a_11279_12268# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3095 a_9888_16532# a_5612_17317# vccd1 vccd1 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3096 a_4698_22020# a_4578_21976# a_3954_21976# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3097 a_3319_21237# a_2500_22020# a_3507_21237# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3098 vccd1 a_3212_11872# a_3108_11916# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3099 a_4348_7909# a_5577_9040# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3100 a_27452_19624# a_27364_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3101 a_7404_9006# a_8300_8648# a_8212_8693# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3102 vccd1 a_15804_7080# a_15716_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3103 a_23196_5512# a_23108_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D108 vssd1 a_2140_17302# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3104 a_7302_10836# a_6470_10260# a_7134_10836# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3105 a_8156_17584# a_9800_18056# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3106 a_10136_13396# a_9076_15704# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3107 vccd1 a_6440_18056# a_1692_18528# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3108 vssd1 a_10808_17662# a_10616_17775# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3109 a_1772_23544# a_3564_23544# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3110 vccd1 a_22748_19624# a_22660_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3111 a_13496_15774# a_14708_18100# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X3112 a_7292_9880# a_7192_9710# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3113 a_7884_24328# a_9519_22020# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X3114 a_20172_18056# a_20084_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3115 a_25884_3511# a_25796_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3116 a_7337_25940# a_6607_25962# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X3117 a_10320_17360# a_11548_13824# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3118 vccd1 a_10036_16532# a_10740_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X3119 vccd1 a_21404_13352# a_21316_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3120 a_20060_7080# a_19972_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3121 vccd1 a_3036_3944# a_2948_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3122 vccd1 a_16140_9783# a_16052_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3123 a_7292_9880# a_7192_9710# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3124 a_19612_16488# a_19524_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3125 vccd1 a_4233_20016# a_4128_20156# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X3126 vccd1 a_16140_6647# a_16052_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3127 vccd1 a_27452_25896# a_27364_25940# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3128 a_9800_18056# a_11628_18056# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X3129 vccd1 a_11548_13824# a_11460_13880# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3130 a_22076_3511# a_21988_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3131 a_13900_8648# a_13812_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3132 a_6383_25940# a_5759_25940# a_6215_25940# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3133 vccd1 a_27452_22760# a_27364_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3134 a_5972_17720# a_5524_17361# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3135 a_16192_25244# a_14471_25571# a_15064_25502# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3136 a_20260_23588# a_19556_23992# vccd1 vccd1 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
D109 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3137 a_26556_7080# a_26468_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3138 vccd1 a_24876_17623# a_24788_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3139 a_7535_11503# a_6635_11000# vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3140 a_10224_24372# a_8492_24328# vccd1 vccd1 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3141 vssd1 a_4481_24757# a_18435_24860# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X3142 a_9856_22875# a_9444_23288# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3143 a_20060_19191# a_19972_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3144 a_10752_12700# a_10604_12967# a_10584_12700# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3145 a_22188_8215# a_22100_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3146 SDAC[2] a_1772_9432# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3147 vccd1 a_17372_14920# a_17284_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3148 vccd1 a_10988_5079# a_10900_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3149 SDAC[1] a_1772_6296# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3150 vccd1 a_17372_11784# a_17284_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3151 a_6531_15357# a_6861_15429# a_6981_14986# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3152 a_13116_3944# a_13028_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3153 SDAC[0] a_1772_3160# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3154 vccd1 a_27900_21192# a_27812_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3155 a_2364_18188# a_2264_18144# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3156 a_3360_8763# a_2948_9176# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3157 vccd1 a_24092_10216# a_24004_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3158 vccd1 a_5612_5079# a_5524_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3159 a_25324_6647# a_25236_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3160 a_16112_20540# a_14000_20856# a_15800_20540# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3161 a_19500_17623# a_19412_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3162 vccd1 a_8568_7930# a_3564_6296# vccd1 pfet_06v0 ad=0.458p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
D110 a_2220_24686# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3163 vccd1 a_27452_16488# a_27364_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D111 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3164 vccd1 a_19357_23336# a_19477_22804# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3165 a_22300_19624# a_22212_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3166 a_3816_15452# a_1604_15448# a_2876_15008# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3167 vccd1 a_17820_13352# a_17732_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3168 vssd1 a_1772_12568# SDAC[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3169 vccd1 a_14908_3944# a_14820_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3170 a_13440_21724# a_13292_21280# a_13272_21724# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3171 vccd1 a_2220_24686# a_17585_20856# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3172 vccd1 a_9920_20096# a_4815_20408# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3173 vccd1 a_10604_25511# a_10500_25560# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3174 a_1996_11000# a_10584_22042# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3175 a_3524_24460# a_3404_24812# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X3176 a_23644_16488# a_23556_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3177 a_9532_3944# a_9444_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3178 a_11525_24164# a_11405_23544# a_10781_23544# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3179 vccd1 a_8752_8648# a_8212_8693# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3180 vccd1 a_23308_18056# a_23220_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D112 a_1692_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3181 a_8156_17584# a_9800_18056# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3182 vccd1 a_14428_23544# a_14272_23992# vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X3183 vssd1 a_1916_17302# a_9572_18884# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3184 vccd1 a_6440_18056# a_1692_18528# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3185 a_19477_23380# a_19357_23336# a_18733_23269# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3186 a_13496_15774# a_14708_18100# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X3187 a_20172_14487# a_20084_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3188 vccd1 a_17372_3511# a_17284_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3189 a_23980_8215# a_23892_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3190 vssd1 a_10584_22042# a_1996_11000# vssd1 nfet_06v0 ad=0.151p pd=1.185u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3191 a_4573_17272# a_2544_19306# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3192 vccd1 a_24092_3944# a_24004_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3193 a_17708_11351# a_17620_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3194 vssd1 a_10732_24328# a_15940_26471# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3195 a_11525_23588# a_11405_23544# a_10781_23544# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3196 a_4573_14136# a_4965_14136# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3197 vccd1 a_10604_12967# a_10500_13016# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3198 a_6635_11000# a_6983_11268# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X3199 vccd1 a_10716_22848# a_10612_22892# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3200 a_6907_23380# a_6431_22804# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3201 vssd1 a_22604_21976# a_22556_22020# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3202 vccd1 a_20732_21192# a_20644_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3203 vccd1 a_4815_20408# a_8736_19363# vccd1 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3204 a_23532_17623# a_23444_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3205 a_20060_3511# a_19972_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3206 vccd1 a_11772_7080# a_11684_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3207 DIGITAL_OUT[0] a_9408_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3208 a_4913_24860# a_2724_24856# a_4041_24812# vccd1 pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X3209 a_10540_5079# a_10452_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3210 a_10901_23588# a_10781_23544# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3211 vccd1 a_21852_13352# a_21764_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3212 a_24540_7080# a_24452_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3213 a_5237_10261# a_4233_10608# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3214 vssd1 a_1772_25112# SC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3215 vccd1 a_17452_20108# a_12860_21976# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3216 vccd1 a_7516_3944# a_7428_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3217 vccd1 a_26668_23895# a_26580_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3218 a_11011_15704# a_11341_15704# a_11461_16302# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3219 a_20172_8215# a_20084_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3220 a_6742_10836# a_6266_10260# a_6470_10260# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3221 a_12650_11828# a_12026_11828# a_12482_11828# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3222 a_15800_25244# a_14872_25615# a_15632_25244# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3223 vssd1 a_10451_23544# a_8456_23632# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3224 a_15568_23992# a_15156_23671# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3225 vccd1 a_26668_20759# a_26580_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3226 a_4578_21976# a_4315_21237# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3227 a_4815_20408# a_9920_20096# vssd1 vssd1 nfet_06v0 ad=0.1248p pd=1u as=0.1248p ps=1u w=0.48u l=0.6u
X3228 a_2588_5512# a_2500_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3229 a_18256_25560# a_17844_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3230 a_25648_25560# a_20652_22424# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3231 a_8548_18884# a_5836_22760# a_9164_18884# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3232 vccd1 a_6719_16532# a_7175_16554# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3233 a_26668_8215# a_26580_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3234 a_6796_25511# a_6488_25560# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3235 vccd1 a_22300_16488# a_22212_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3236 vssd1 a_11961_25200# a_11856_25244# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3237 vccd1 a_5836_22760# a_9076_15704# vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3238 vccd1 a_13048_16576# a_12856_16620# vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3239 vccd1 a_4578_21976# a_4698_22596# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3240 a_3823_18885# a_3703_18840# a_3228_17317# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3241 vccd1 a_3036_5079# a_2948_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3242 vccd1 a_16140_8648# a_16052_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3243 a_5472_9180# a_2948_9176# a_5160_9180# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3244 a_4128_23292# a_1604_23288# a_3816_23292# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3245 a_4128_18588# a_2016_18171# a_3816_18588# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3246 a_10408_22892# a_9856_22875# a_10204_22892# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3247 a_12911_19756# a_11787_20027# vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3248 vccd1 a_26668_14487# a_26580_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3249 vccd1 a_24876_9783# a_24788_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3250 a_4716_25204# a_11961_25200# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3251 a_4128_20156# a_1604_20152# a_3816_20156# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3252 vccd1 a_5544_7584# a_3564_12568# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3253 a_7646_19438# a_7190_18884# a_7414_18884# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3254 a_1692_18528# a_6440_18056# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3255 vccd1 a_24876_6647# a_24788_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3256 vccd1 a_26668_11351# a_26580_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3257 vccd1 a_6796_25511# a_6692_25560# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3258 a_2876_22848# a_2568_22892# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3259 vccd1 a_15468_11351# a_15380_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3260 a_5573_11829# a_4569_12176# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3261 vssd1 a_5627_23544# a_5539_23589# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3262 vssd1 a_1772_12568# SDAC[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3263 a_20112_24860# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3264 a_9295_22596# a_8671_22020# a_9127_22596# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3265 a_2876_19712# a_2568_19756# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3266 a_11628_18056# a_13496_17337# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3267 vssd1 a_9123_17317# a_10900_14964# vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3268 vccd1 a_2668_9132# a_2264_15008# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3269 SDAC[5] a_1772_20408# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3270 a_13572_13016# a_8435_13397# vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X3271 a_5559_11448# a_5831_11000# a_5132_7564# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3272 vssd1 a_13497_14964# a_14176_17020# vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3273 vssd1 a_5817_24800# a_5769_24856# vssd1 nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X3274 a_19428_23588# a_19308_23544# vssd1 vssd1 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3275 a_25660_5512# a_25572_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3276 a_2672_21782# a_1916_22021# vssd1 vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X3277 vccd1 a_27116_17623# a_27028_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3278 a_21292_6647# a_21204_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3279 a_3072_10564# a_9744_8392# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3280 vccd1 a_4731_20872# a_10104_22848# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3281 a_9846_20152# a_5836_22760# a_9652_20152# vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X3282 vccd1 a_23756_18056# a_23668_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3283 a_9644_5079# a_9556_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3284 a_6839_25962# a_6383_25940# a_6607_25962# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3285 a_6859_20452# a_6383_21028# a_6607_20452# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3286 vccd1 a_5019_20408# a_9076_15704# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3287 vccd1 a_21740_19191# a_21652_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3288 vccd1 a_20508_10216# a_20420_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3289 a_8352_23676# a_6631_24003# a_7224_23934# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3290 a_12158_11784# a_11961_12656# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3291 vccd1 a_8153_25200# a_8048_25244# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X3292 a_1812_17353# a_2140_17302# a_2016_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3293 vccd1 a_10876_3944# a_10788_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3294 COMP_CLK a_2444_26249# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3295 a_8736_19363# a_4815_20408# vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3296 a_27004_18056# a_26916_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3297 a_15351_24394# a_14895_24372# a_15119_24394# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3298 a_25324_23895# a_25236_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3299 a_23868_21192# a_23780_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3300 a_27004_14920# a_26916_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3301 a_4693_11620# a_4573_11000# a_3949_11000# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3302 a_6488_25560# a_5936_25560# a_6284_25560# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3303 a_1772_11000# a_5831_11000# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3304 vssd1 a_18403_21629# a_17452_20108# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3305 a_19724_12919# a_19636_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3306 a_4964_9880# a_4516_9521# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3307 a_11669_24856# a_4631_20408# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3308 a_2444_18840# a_8144_19288# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3309 vccd1 a_23644_8648# a_23556_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3310 a_8756_18884# a_5836_22760# a_8548_18884# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3311 a_23980_17623# a_23892_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3312 a_24540_3511# a_24452_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3313 vssd1 a_9612_15704# a_8972_15749# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3314 vccd1 a_23644_5512# a_23556_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3315 a_9744_8392# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3316 vccd1 a_17372_8648# a_17284_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3317 a_3564_6296# a_8568_7930# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X3318 a_20260_23588# a_19556_23992# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3319 vccd1 a_1916_17302# a_9532_19624# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3320 vccd1 a_17372_5512# a_17284_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3321 vccd1 a_23420_22327# a_23332_22424# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3322 a_13292_21280# a_12984_21324# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3323 a_7784_9564# a_6944_9880# a_7496_9880# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
D113 a_5940_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3324 a_18380_8215# a_18292_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3325 vccd1 a_5020_15796# a_9532_13685# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3326 a_4380_5079# a_4292_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3327 a_25212_7080# a_25124_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3328 a_25648_25560# a_20652_22424# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3329 vssd1 a_9920_20096# a_4815_20408# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
X3330 vccd1 a_3484_3944# a_3396_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3331 vccd1 a_3816_13884# a_4233_13744# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X3332 vccd1 a_1692_17302# a_14986_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3333 vssd1 a_3072_10564# a_3360_12316# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3334 a_27228_3511# a_27140_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3335 a_18268_19191# a_18180_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3336 a_8624_14602# a_7281_7142# a_8644_14181# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3337 vssd1 a_2444_24328# a_7572_24856# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3338 vssd1 a_3072_10564# a_4368_9180# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3339 vccd1 CLK a_13496_17337# vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3340 a_3932_7080# a_3844_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3341 a_4180_18884# a_4492_18840# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3342 a_11909_9476# a_11789_9432# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3343 a_1772_20408# a_3564_20408# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3344 a_10808_17662# a_10320_17360# a_11068_17720# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3345 a_5948_3511# a_5860_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3346 vccd1 a_4264_17020# a_4681_16880# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X3347 a_4152_12316# a_1940_12312# a_3212_11872# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3348 a_13564_3944# a_13476_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3349 a_12152_10304# a_11559_10304# a_12888_10748# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3350 a_5076_23992# a_4628_23633# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3351 vccd1 a_27564_17623# a_27476_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3352 a_25772_6647# a_25684_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D114 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3353 vccd1 a_22476_25511# a_22372_25560# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3354 vssd1 a_9800_18056# a_8156_17584# vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3355 vssd1 a_13496_17337# a_11628_18056# vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3356 vccd1 a_17932_14487# a_17844_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3357 a_23196_7080# a_23108_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3358 a_3682_22020# a_3542_22242# a_2918_21976# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3359 vccd1 a_19276_9783# a_19188_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3360 DIGITAL_OUT[5] a_24640_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3361 a_4913_24860# a_3136_24443# a_4041_24812# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X3362 a_27900_22760# a_27812_22804# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3363 vccd1 a_19276_6647# a_19188_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3364 vssd1 a_13216_25940# DIGITAL_OUT[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3365 vssd1 a_4731_20872# a_20299_21720# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3366 vssd1 a_14708_18100# a_15456_19368# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3367 vccd1 a_20956_10216# a_20868_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3368 vssd1 a_21392_25940# DIGITAL_OUT[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3369 vccd1 a_12262_23544# a_5940_6390# vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3370 vssd1 a_7190_18884# a_7666_18884# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3371 a_11459_11000# a_11789_11000# a_11909_11044# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3372 COMP_CLK a_2444_26249# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3373 vssd1 a_13776_18100# a_14708_18100# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3374 a_27452_18056# a_27364_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3375 a_25772_23895# a_25684_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3376 a_27452_14920# a_27364_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3377 vccd1 a_5836_22760# a_2444_24328# vccd1 pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3378 vccd1 a_5237_18101# a_5530_18884# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3379 vccd1 a_14348_8215# a_14260_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3380 vccd1 a_16812_16055# a_16724_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3381 a_9980_3944# a_9892_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3382 vccd1 a_2444_24328# a_1996_24328# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3383 vccd1 a_13252_22804# a_9900_24756# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3384 vssd1 a_12108_21664# a_15156_23671# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3385 vccd1 a_3542_22242# a_3642_22596# vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3386 a_12337_25244# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3387 vssd1 a_13077_22805# a_15940_22065# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3388 a_4684_7564# a_5831_12568# a_5767_12613# vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3389 vccd1 a_8748_5079# a_8660_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3390 a_8764_15749# a_9123_17317# a_9176_16177# vccd1 pfet_06v0 ad=0.4012p pd=1.85u as=0.58035p ps=2.155u w=1.095u l=0.5u
X3391 a_22168_25560# a_21616_25560# a_21964_25560# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3392 vccd1 a_14649_21584# a_5836_22760# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3393 vccd1 a_15456_19368# a_12108_21664# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3394 vccd1 a_14392_14181# a_8335_13352# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3395 a_6172_3944# a_6084_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3396 vccd1 a_5237_10261# a_5642_10260# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3397 a_16744_22042# a_16388_22424# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.151p ps=1.185u w=0.36u l=0.6u
X3398 a_18403_21629# a_18733_21701# a_18853_21258# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3399 vccd1 a_20396_17623# a_20308_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3400 vccd1 a_8437_10291# a_8247_13397# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3401 a_26108_21192# a_26020_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D115 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3402 vccd1 a_24092_14920# a_24004_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3403 vccd1 a_15392_13824# a_8519_13836# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3404 vccd1 a_13292_21280# a_13188_21324# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3405 vccd1 a_7259_24800# a_2444_24328# vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.52205p ps=2.045u w=0.985u l=0.5u
X3406 vccd1 a_24092_11784# a_24004_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3407 a_7511_11850# a_7055_11828# a_7279_11850# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3408 a_7337_20856# a_6607_20452# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
D116 vssd1 a_5940_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3409 a_4684_7564# a_4964_9880# a_5559_13016# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3410 vccd1 a_7964_3944# a_7876_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3411 a_25324_8215# a_25236_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3412 vccd1 a_23420_21192# a_23332_21236# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3413 a_3816_20156# a_1604_20152# a_2876_19712# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3414 a_26220_17623# a_26132_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3415 vssd1 a_7302_14180# a_7778_14180# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3416 a_7988_3608# a_7540_3249# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3417 vccd1 a_13116_7080# a_13028_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3418 vccd1 a_23532_9783# a_23444_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3419 vssd1 a_5940_6390# a_5600_18101# vssd1 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X3420 vccd1 a_24540_13352# a_24452_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3421 vssd1 a_4481_24757# a_13440_21724# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3422 vccd1 a_23532_6647# a_23444_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3423 a_13920_23992# a_13820_23544# vccd1 vccd1 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3424 vccd1 a_27900_19624# a_27812_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3425 a_6383_21028# a_5759_20452# a_6235_20452# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3426 a_24428_20759# a_24340_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3427 a_2812_16620# a_2712_16576# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3428 vccd1 a_1772_9432# SDAC[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3429 a_26108_11784# a_26020_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3430 vccd1 a_23644_23291# a_23556_23335# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X3431 vccd1 a_3484_5079# a_3396_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3432 vccd1 a_1772_6296# SDAC[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3433 a_10192_8692# a_7988_3608# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3434 a_10684_24856# a_9900_24756# a_10372_24372# vssd1 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3435 a_7032_24047# a_6736_23632# a_5975_23812# vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3436 a_7744_11088# a_1692_10688# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3437 a_11909_11598# a_11789_11000# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X3438 a_4569_12176# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X3439 a_8435_13397# a_8335_13352# a_8247_13397# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3440 vccd1 a_1772_3160# SDAC[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3441 a_22300_14920# a_22212_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3442 a_4945_12316# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3443 vccd1 a_28012_5079# a_27924_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3444 DIGITAL_OUT[5] a_24640_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3445 a_12108_21664# a_15456_19368# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3446 a_20508_3944# a_20420_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3447 a_8444_24856# a_2444_24328# a_8132_24372# vssd1 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3448 a_17708_16055# a_17620_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3449 a_8300_5079# a_8212_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3450 vssd1 a_13216_25940# DIGITAL_OUT[1] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3451 vssd1 a_21392_25940# DIGITAL_OUT[4] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3452 a_24428_14487# a_24340_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3453 a_9537_9564# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3454 vccd1 a_9295_22596# a_9751_22574# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3455 a_5139_21292# a_4403_21582# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3276p ps=1.62u w=0.78u l=0.5u
X3456 vccd1 a_14860_20807# a_14756_20856# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3457 a_4233_13744# a_3816_13884# a_4609_13884# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3458 vssd1 a_9076_15704# a_11032_13880# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3459 a_24428_11351# a_24340_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3460 a_8548_18884# a_4815_20408# a_10884_18884# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3461 vccd1 a_18828_8215# a_18740_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3462 a_3072_10564# a_9744_8392# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3463 a_4233_10608# a_3816_10748# a_4609_10748# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3464 vccd1 a_18156_11351# a_18068_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D117 a_2140_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3465 vccd1 a_17947_24328# a_17859_24373# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3466 a_10240_16532# a_9476_17016# a_10036_16532# vccd1 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3467 a_4716_18840# a_4233_15312# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3468 vccd1 a_1772_25112# SC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3469 a_14708_18100# a_13776_18100# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3470 a_3708_8780# a_3608_8736# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3471 a_10676_16152# a_10228_15793# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3472 a_12220_13484# a_10808_13880# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3473 a_13900_9783# a_13812_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3474 a_2444_24328# a_5836_22760# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3475 vccd1 a_22300_8648# a_22212_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3476 a_19477_18676# a_19357_18632# a_18733_18565# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3477 vccd1 a_3072_10564# a_9211_17272# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X3478 vssd1 CLK a_13496_17337# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3479 vccd1 a_22300_5512# a_22212_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3480 a_27004_5512# a_26916_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3481 vccd1 a_17036_12919# a_16948_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3482 vssd1 a_5940_6390# a_6299_7608# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3483 a_2588_7080# a_2500_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3484 vssd1 a_2668_9132# a_2264_15008# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3485 vccd1 a_22188_20759# a_22100_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3486 vccd1 a_15456_19368# a_12108_21664# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3487 a_18853_18675# a_18733_18565# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3488 vssd1 a_5836_22760# a_11676_20452# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X3489 a_9180_14609# a_6388_6390# a_8868_14609# vccd1 pfet_06v0 ad=0.2847p pd=1.615u as=0.58035p ps=2.155u w=1.095u l=0.5u
X3490 a_6175_12613# a_3703_18840# a_4684_7564# vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3491 vssd1 a_10159_10700# a_10095_10744# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3492 a_14552_20856# a_13588_20535# a_14348_20856# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3493 a_28012_23895# a_27924_23992# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3494 a_26556_21192# a_26468_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3495 a_8736_19363# a_10452_18840# a_10378_18884# vssd1 nfet_06v0 ad=0.4161p pd=1.905u as=0.1517p ps=1.19u w=0.82u l=0.6u
X3496 a_6172_9432# a_5831_12568# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3497 a_5724_5512# a_5636_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3498 a_14552_20856# a_14000_20856# a_14348_20856# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3499 vccd1 a_1772_15704# SDAC[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3500 a_11548_13824# a_13496_15774# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3501 vccd1 a_6060_23118# a_3404_24812# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3502 vccd1 a_13496_15774# a_11548_13824# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3503 vccd1 a_1772_12568# SDAC[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3504 a_6590_19460# a_6154_19460# a_6358_19378# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3505 vccd1 a_5237_19669# a_5759_20452# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3506 vccd1 a_2140_3944# a_2052_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3507 vccd1 a_22188_14487# a_22100_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3508 a_12432_21307# a_12020_21720# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3509 vccd1 a_21392_25940# DIGITAL_OUT[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3510 vccd1 a_22188_11351# a_22100_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3511 a_21180_3511# a_21092_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3512 vccd1 a_20776_24766# a_20672_24860# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3513 a_6702_14756# a_6266_14756# a_6470_14674# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3514 a_3981_24460# a_2724_24856# a_3728_24460# vccd1 pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X3515 a_25660_7080# a_25572_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3516 a_24876_20759# a_24788_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3517 a_4128_18588# a_1604_18584# a_3816_18588# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3518 a_4693_14180# a_4573_14136# a_3949_14136# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3519 a_21292_8215# a_21204_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3520 SDAC[2] a_1772_9432# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3521 a_26556_11784# a_26468_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3522 a_4604_6647# a_4516_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3523 a_15356_11784# a_15268_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3524 vccd1 a_20508_14920# a_20420_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3525 a_27676_3511# a_27588_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3526 SDAC[1] a_1772_6296# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3527 vccd1 a_19612_10216# a_19524_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3528 a_4693_11044# a_4573_11000# a_3949_11000# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3529 a_11011_15704# a_11341_15704# a_11461_15748# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3530 a_4604_3511# a_4516_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3531 a_24640_25940# a_24004_22804# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3532 a_2876_18144# a_2568_18188# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3533 a_12220_3944# a_12132_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3534 SDAC[0] a_1772_3160# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3535 vccd1 a_20508_11784# a_20420_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3536 vccd1 a_5084_25560# a_13216_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3537 a_13188_21324# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X3538 a_8232_11390# a_7744_11088# a_8492_11448# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3539 a_24004_22804# a_23556_23335# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3540 SDAC[4] a_1772_15704# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3541 a_5544_7584# a_5573_11829# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X3542 vccd1 a_2444_24328# a_7852_9006# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3543 a_12984_21324# a_12020_21720# a_12780_21324# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3544 a_1812_17353# a_1692_17302# vssd1 vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X3545 a_24876_14487# a_24788_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3546 a_6523_20243# a_6047_19668# a_6271_19690# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3547 a_18716_3944# a_18628_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3548 a_24876_11351# a_24788_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3549 a_13776_18100# a_11628_18056# vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3550 vssd1 a_1812_17353# a_5412_15495# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3551 a_9800_14181# a_8624_14602# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X3552 a_14348_5079# a_14260_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3553 vccd1 a_3564_23544# a_1772_23544# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3554 a_9800_18056# a_11628_18056# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X3555 a_8009_11828# a_7279_11850# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X3556 vssd1 a_14576_25200# a_14471_25571# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3557 a_19544_24416# a_19056_24816# a_19804_24460# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3558 vccd1 a_13900_12568# a_12581_14136# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3559 vccd1 a_3564_20408# a_1772_20408# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3560 vccd1 a_8156_17584# a_6440_18056# vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
D118 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3561 DIGITAL_OUT[3] a_18256_25560# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3562 vccd1 a_16773_18528# a_9612_15704# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3563 COMP_CLK a_2444_26249# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3564 a_7736_25244# a_5524_25239# a_6796_25511# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3565 a_5685_16533# a_4681_16880# vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3566 a_10662_20152# a_9920_20096# a_10468_20152# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X3567 vssd1 a_3072_10564# a_3024_13884# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3568 vccd1 a_17484_12919# a_17396_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3569 vccd1 a_14796_8215# a_14708_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3570 vccd1 a_22188_9783# a_22100_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3571 SC a_1772_25112# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3572 a_5895_21372# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.1521p pd=1.105u as=0.4149p ps=2.65u w=0.585u l=0.5u
X3573 vssd1 a_1692_10688# a_9332_12695# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3574 vccd1 a_7404_5079# a_7316_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3575 a_27116_6647# a_27028_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3576 vccd1 a_22188_6647# a_22100_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3577 vssd1 a_9744_8392# a_3072_10564# vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3578 a_7055_11828# a_6431_11828# a_6887_11828# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3579 vssd1 a_3072_10564# a_3024_10748# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3580 a_24209_25244# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3581 a_16388_22424# a_15940_22065# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3582 vccd1 a_23644_10216# a_23556_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3583 a_9540_12268# a_6388_6390# vssd1 vssd1 nfet_06v0 ad=0.14p pd=1.1u as=0.224p ps=1.52u w=0.4u l=0.6u
X3584 a_11960_10348# a_11559_10304# a_10903_10216# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3585 a_1692_18528# a_6440_18056# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3586 a_13672_13884# a_11872_13467# a_12732_13440# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3587 a_5160_9180# a_2948_9176# a_4220_8736# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3588 vccd1 a_19500_16055# a_19412_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3589 a_5831_12568# a_7526_14180# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X3590 vssd1 a_7744_11088# a_7639_11459# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3591 a_2220_14136# a_4492_18840# a_4388_19288# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3592 a_23221_24394# a_23101_24837# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X3593 a_14392_14181# a_5972_17720# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X3594 vccd1 a_6620_3944# a_6532_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3595 vssd1 a_1772_23544# SDAC[6] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3596 vccd1 a_6736_23632# a_6631_24003# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3597 a_7485_13928# a_5573_11829# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3598 a_8420_9176# a_8300_8648# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3599 a_21404_11784# a_21316_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3600 a_16217_20496# a_15800_20540# a_16593_20540# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3601 SDAC[4] a_1772_15704# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3602 vssd1 a_13496_15774# a_11548_13824# vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3603 vccd1 a_21392_25940# DIGITAL_OUT[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3604 a_14576_25200# a_12108_21664# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3605 EOC a_25648_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3606 vssd1 a_14895_24372# a_15371_24947# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3607 vssd1 a_12650_11828# a_13126_12404# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3608 SDAC[3] a_1772_12568# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3609 vccd1 a_25436_3511# a_25348_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3610 a_6944_25244# a_6796_25511# a_6776_25244# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3611 vssd1 a_9211_17272# a_9123_17317# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3612 a_1692_5512# a_1604_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D119 vssd1 a_2444_24328# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3613 vccd1 a_7485_13928# a_7605_13396# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3614 a_3564_6296# a_8568_7930# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3615 a_2164_21236# a_1716_21767# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3616 vccd1 a_3619_17272# a_2264_18144# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3617 vccd1 a_19164_3511# a_19076_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3618 vccd1 a_14708_18100# a_15456_19368# vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3619 a_25772_8215# a_25684_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3620 a_5612_23118# a_7259_24800# a_16709_21720# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3621 vccd1 a_2444_24328# a_13900_12568# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3622 vccd1 a_20956_14920# a_20868_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3623 vccd1 a_23084_17623# a_22996_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3624 a_6531_13789# a_6861_13861# a_6981_13971# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3625 vccd1 a_2140_5079# a_2052_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3626 a_13467_25112# a_13815_25380# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X3627 a_16700_3944# a_16612_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3628 vccd1 a_13564_7080# a_13476_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3629 vccd1 a_20956_11784# a_20868_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3630 a_10616_17775# a_10215_17731# a_9559_17540# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3631 vccd1 a_23980_9783# a_23892_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3632 a_12332_5079# a_12244_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3633 a_1772_15704# a_3564_15704# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3634 vccd1 a_23980_6647# a_23892_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3635 vccd1 a_27197_24904# a_27317_24372# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3636 vccd1 a_1772_9432# SDAC[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3637 vccd1 a_10428_11351# a_10340_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3638 a_2444_24328# a_7259_24800# a_9560_20452# vssd1 nfet_06v0 ad=0.4161p pd=1.905u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3639 a_13497_14964# a_12767_14986# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X3640 a_10320_17360# a_11548_13824# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3641 vccd1 a_23532_16055# a_23444_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3642 a_2904_11916# a_2352_11899# a_2700_11916# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3643 vccd1 a_1772_6296# SDAC[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3644 a_8849_10744# a_2220_24686# a_8645_10744# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.1722p ps=1.24u w=0.82u l=0.6u
X3645 a_17820_11784# a_17732_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3646 vccd1 a_1772_3160# SDAC[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3647 vccd1 a_23532_12919# a_23444_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3648 a_18828_5079# a_18740_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3649 a_10555_21267# a_9900_13396# vccd1 vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3650 vccd1 a_20172_9783# a_20084_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3651 a_6527_24047# a_5627_23544# vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3652 a_27116_20759# a_27028_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3653 vssd1 a_5880_12288# a_1692_18885# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X3654 vccd1 a_8156_17584# a_6440_18056# vccd1 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3655 vccd1 a_20172_6647# a_20084_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3656 a_20956_3944# a_20868_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3657 vssd1 a_18256_25560# DIGITAL_OUT[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3658 a_5472_9180# a_3360_8763# a_5160_9180# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3659 a_5139_21292# a_3072_10564# a_5159_21720# vssd1 nfet_06v0 ad=0.3123p pd=2.38u as=48.6f ps=0.645u w=0.405u l=0.6u
X3660 a_4233_23152# a_3816_23292# a_4609_23292# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3661 vccd1 a_4760_12613# a_4672_12657# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3662 vccd1 a_26668_9783# a_26580_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3663 a_1772_25112# a_3564_25112# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3664 a_4233_20016# a_3816_20156# a_4609_20156# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3665 vccd1 a_26668_6647# a_26580_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3666 a_7628_5512# a_7540_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3667 a_11872_13467# a_11460_13880# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3668 a_1692_10688# a_6328_17342# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3669 a_3472_17020# a_3324_16576# a_3304_17020# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3670 a_27116_14487# a_27028_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3671 a_3319_21237# a_3999_21676# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3672 vccd1 a_7055_11828# a_7511_11850# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3673 a_23416_25244# a_21204_25239# a_22476_25511# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3674 a_27116_11351# a_27028_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3675 vssd1 a_10372_24372# a_11076_24372# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3676 a_8225_14965# a_5972_17720# a_8617_15448# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3677 vccd1 a_23420_3511# a_23332_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3678 a_27452_5512# a_27364_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3679 a_3004_21664# a_5836_22760# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X3680 a_10555_21267# a_2220_24686# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X3681 vssd1 a_9532_13685# a_9444_13880# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3682 a_23084_6647# a_22996_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D120 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3683 a_13120_20112# a_12108_21664# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3684 a_13048_16576# a_12455_16576# a_13784_17020# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3685 a_4368_9180# a_4220_8736# a_4200_9180# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3686 a_10348_15448# a_9900_13396# a_9532_19624# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3687 a_21852_11784# a_21764_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3688 a_15324_25560# a_14872_25615# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X3689 a_2568_13484# a_1604_13880# a_2364_13484# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3690 a_16520_20128# COMP_OUT vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X3691 a_1772_15704# a_3564_15704# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3692 a_2568_10348# a_1604_10744# a_2364_10348# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3693 vccd1 a_20060_13352# a_19972_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3694 a_1772_12568# a_3564_12568# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3695 vccd1 a_12668_3944# a_12580_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3696 vccd1 a_13832_15424# a_5612_17317# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3697 a_14348_8648# a_14260_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3698 vccd1 a_26108_18056# a_26020_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3699 DIGITAL_OUT[4] a_21392_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3700 a_7531_23379# a_7055_22804# a_7279_22826# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3701 a_6981_13418# a_6861_13861# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X3702 vccd1 a_6328_17342# a_1692_10688# vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3703 a_12308_22020# a_9532_19624# a_12100_22020# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3704 a_24428_19191# a_24340_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3705 vssd1 a_1772_9432# SDAC[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3706 a_22624_25244# a_22476_25511# a_22456_25244# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3707 a_26332_3511# a_26244_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3708 a_3038_22020# a_2918_21976# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3709 a_24428_16055# a_24340_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3710 a_8225_14965# a_4492_18840# vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3711 vssd1 a_8721_14920# a_10136_13396# vssd1 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3712 a_21740_12919# a_21652_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3713 vccd1 a_19164_8648# a_19076_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3714 a_8437_10291# a_2220_24686# vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3715 a_6383_25940# a_5759_25940# a_6235_26516# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3716 a_19164_13352# a_19076_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3717 vssd1 a_3564_23544# a_1772_23544# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3718 vccd1 a_19164_5512# a_19076_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3719 a_12413_9432# a_8752_8648# vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3720 vccd1 a_26668_19191# a_26580_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3721 a_12220_13484# a_10808_13880# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3722 vccd1 a_20508_7080# a_20420_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3723 a_19164_10216# a_19076_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3724 a_13086_11828# a_12650_11828# a_12854_11828# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3725 vccd1 a_23980_16055# a_23892_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3726 a_1872_11466# a_1772_11000# vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3727 a_12308_22424# a_9532_19624# vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3728 vccd1 a_6547_11045# a_6543_12612# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3729 vccd1 a_23980_12919# a_23892_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3730 a_22096_22424# a_17859_24373# vccd1 vccd1 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3731 vccd1 a_7302_14180# a_7758_14734# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3732 a_27564_20759# a_27476_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3733 a_4481_24757# a_10192_8692# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3734 a_7778_10835# a_7302_10836# a_7526_10282# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3735 a_27004_7080# a_26916_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3736 SC a_1772_25112# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3737 vssd1 a_5795_21280# a_5547_21551# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3738 vccd1 a_4481_24757# a_13308_16620# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3739 vccd1 a_5276_3944# a_5188_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3740 vccd1 a_18380_9783# a_18292_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3741 vccd1 a_8721_14920# a_10324_13396# vccd1 pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
X3742 SDAC[2] a_1772_9432# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3743 vccd1 a_11436_5079# a_11348_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3744 vccd1 a_18380_6647# a_18292_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3745 vssd1 a_17947_24328# a_17859_24373# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3746 a_24005_24142# a_23885_23544# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X3747 vssd1 a_4578_21976# a_4698_22020# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3748 SDAC[1] a_1772_6296# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3749 vssd1 a_6440_18056# a_1692_18528# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3750 vssd1 a_9920_20096# a_4815_20408# vssd1 nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3751 SDAC[0] a_1772_3160# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3752 a_22412_18056# a_22324_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3753 a_14796_5079# a_14708_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3754 a_9056_9564# a_6944_9880# a_8744_9564# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3755 a_7154_10260# a_6470_10260# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X3756 vccd1 a_5627_23544# a_5539_23589# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3757 vssd1 a_5237_10261# a_5642_10260# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X3758 a_18312_22021# a_2276_22424# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X3759 vccd1 a_13452_8215# a_13364_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D121 vssd1 a_5940_6390# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3760 a_15288_22021# a_12308_22020# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X3761 a_1692_10688# a_6328_17342# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3762 a_27564_14487# a_27476_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D122 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3763 a_22076_21192# a_21988_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3764 a_8144_19288# a_7414_18884# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X3765 vccd1 CLK a_13496_17337# vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3766 vssd1 a_12560_16976# a_12455_16576# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3767 a_27564_11351# a_27476_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3768 a_15356_3944# a_15268_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3769 a_16364_11351# a_16276_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3770 a_4069_17316# a_3949_17272# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3771 vssd1 a_6328_17342# a_1692_10688# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
D123 a_1804_21723# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3772 a_23196_13352# a_23108_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3773 vssd1 a_3072_10564# a_3024_23292# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3774 vccd1 a_7852_5079# a_7764_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3775 a_27564_6647# a_27476_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3776 a_23196_10216# a_23108_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3777 a_19760_23992# a_18996_23588# a_19556_23992# vccd1 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3778 a_13653_24372# a_13533_24904# a_12909_24837# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3779 vssd1 a_19544_24416# a_19352_24460# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3780 vssd1 a_3072_10564# a_3024_20156# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3781 a_19357_23336# a_10732_24328# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3782 vssd1 a_3619_17272# a_2264_18144# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3783 a_10428_5512# a_10340_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3784 SDAC[3] a_1772_12568# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3785 vssd1 a_13496_17337# a_11628_18056# vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3786 a_11292_21192# a_11324_19624# vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3787 vccd1 a_19612_14920# a_19524_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3788 a_2464_16603# a_2052_17016# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3789 a_14176_17020# a_12560_16976# a_13048_16576# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3790 vccd1 a_19612_11784# a_19524_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3791 vccd1 a_10584_22042# a_1996_11000# vccd1 pfet_06v0 ad=0.458p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3792 a_20396_20759# a_20308_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D124 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3793 a_12152_10304# a_11664_10704# a_12412_10348# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3794 vccd1 a_26556_18056# a_26468_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3795 a_25212_13352# a_25124_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3796 a_8744_9564# a_6944_9880# a_7804_9831# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
D125 a_4481_24757# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3797 a_12999_14986# a_12543_14964# a_12767_14986# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3798 vccd1 a_4631_20408# a_11636_21236# vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3799 vssd1 a_7001_19668# a_2264_22848# vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3800 vccd1 a_9744_8392# a_3072_10564# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3801 a_25212_10216# a_25124_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3802 a_17680_23676# a_15156_23671# a_17368_23676# vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3803 vccd1 a_15848_20128# a_3564_20408# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3804 a_24876_19191# a_24788_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3805 a_7496_9880# a_6532_9559# a_7292_9880# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3806 a_24876_16055# a_24788_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3807 vssd1 a_3072_10564# a_10752_12700# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3808 vccd1 a_25884_3511# a_25796_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3809 vccd1 a_12220_7080# a_12132_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3810 a_2276_22424# a_1828_22065# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3811 a_6839_21006# a_6383_21028# a_6607_20452# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3812 a_3324_16576# a_3016_16620# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3813 a_12712_13884# a_11872_13467# a_12424_13484# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3814 a_8583_20856# a_9263_20408# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3815 a_20396_11351# a_20308_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3816 vccd1 a_13608_19712# a_13416_19756# vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3817 a_5953_9180# a_3072_10564# vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3818 a_16588_10216# a_16500_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3819 vccd1 a_18716_7080# a_18628_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3820 a_2588_8215# a_2500_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3821 vccd1 a_26108_8648# a_26020_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3822 SDAC[2] a_1772_9432# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3823 a_22948_22020# a_22244_22424# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3824 vccd1 a_26108_5512# a_26020_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3825 vccd1 a_22076_3511# a_21988_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3826 vccd1 a_9408_25940# DIGITAL_OUT[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3827 vccd1 a_20652_22424# a_25648_25560# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3828 a_6551_16532# a_6095_16532# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3829 a_12780_5079# a_12692_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3830 a_3036_5512# a_2948_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3831 a_7484_23992# a_7032_24047# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X3832 vccd1 a_19648_21976# a_3564_25112# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3833 a_1772_25112# a_3564_25112# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3834 vssd1 a_4403_21582# a_4315_21237# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3835 vccd1 a_12560_16976# a_12455_16576# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3836 vccd1 a_10808_17662# a_10616_17775# vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3837 vccd1 a_23644_14920# a_23556_14964# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3838 a_27116_8215# a_27028_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3839 a_21392_25940# a_20196_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3840 vssd1 a_1692_18528# a_5524_25239# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
D126 a_5940_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3841 vccd1 a_23644_11784# a_23556_11828# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3842 vssd1 a_6440_18056# a_1692_18528# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3843 a_22860_18056# a_22772_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3844 vccd1 a_4828_5512# a_4740_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3845 vccd1 a_1692_10688# a_1604_10744# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3846 a_5795_21280# a_1692_18528# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3847 vccd1 a_13776_18100# a_14708_18100# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3848 vccd1 a_25324_9783# a_25236_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3849 vccd1 a_17932_8215# a_17844_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3850 a_23868_22327# a_23780_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3851 vccd1 a_25324_6647# a_25236_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3852 vccd1 a_2444_24328# a_7572_24856# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3853 a_5559_11448# a_6239_11000# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3854 vccd1 a_26220_16055# a_26132_16152# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3855 vssd1 a_17221_20453# a_20196_22112# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3856 a_22771_24765# a_23101_24837# a_23221_24394# vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3857 vccd1 a_26220_12919# a_26132_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3858 vssd1 a_19357_23336# a_19477_23380# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3859 vssd1 a_7988_19668# a_11348_22065# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3860 a_18380_12919# a_18292_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3861 a_14162_12403# a_13686_12404# a_13910_11850# vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3862 vccd1 a_17024_25940# DIGITAL_OUT[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D127 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3863 vccd1 a_7736_25244# a_8153_25200# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X3864 a_1692_7080# a_1604_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3865 a_14908_5512# a_14820_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3866 a_7055_22804# a_6431_22804# a_6907_23380# vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3867 a_7511_22826# a_7055_22804# a_7279_22826# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3868 vssd1 a_1692_18885# a_1604_18929# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3869 vssd1 a_1916_17302# a_4180_18884# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3870 a_12108_21664# a_15456_19368# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3871 vccd1 a_27900_8648# a_27812_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3872 vccd1 a_5940_6390# a_1772_14136# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3873 vccd1 a_12650_11828# a_13086_11828# vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3874 a_10604_12967# a_10296_13016# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X3875 vccd1 a_11324_3944# a_11236_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3876 vccd1 a_27900_5512# a_27812_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3877 a_13004_8648# a_12916_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3878 a_3136_24443# a_2724_24856# vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3879 a_10584_22042# a_9444_19668# vccd1 vccd1 pfet_06v0 ad=0.4488p pd=2.92u as=0.458p ps=2.02u w=1.02u l=0.5u
X3880 a_6328_17342# a_8156_17584# vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X3881 a_25660_13352# a_25572_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3882 a_4041_24812# a_4481_24757# a_4385_24860# vssd1 nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X3883 vccd1 a_5940_6390# a_5412_18101# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3884 vccd1 a_18268_13352# a_18180_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3885 a_13488_11000# a_8927_13836# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X3886 a_25660_10216# a_25572_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3887 a_2568_22892# a_1604_23288# a_2364_22892# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3888 vccd1 a_15800_20540# a_16217_20496# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X3889 a_9652_20152# a_9532_19624# vssd1 vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3890 vccd1 a_20172_14487# a_20084_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3891 vssd1 a_24640_25940# DIGITAL_OUT[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3892 vccd1 a_24092_19624# a_24004_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D128 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3893 vccd1 a_17708_11351# a_17620_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3894 a_11856_25244# a_9744_25560# a_11544_25244# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3895 a_2568_19756# a_1604_20152# a_2364_19756# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3896 a_15456_19368# a_14708_18100# vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3897 a_14380_23588# a_9900_24756# a_14068_23992# vssd1 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3898 vssd1 a_2444_26249# COMP_CLK vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3899 vssd1 a_14428_23544# a_17396_25201# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3900 vccd1 a_22604_21976# a_22448_22424# vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X3901 a_14708_18100# a_13776_18100# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X3902 vccd1 a_16700_7080# a_16612_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3903 a_14796_8648# a_14708_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3904 vccd1 a_13120_20112# a_13015_19712# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3905 vccd1 a_20060_3511# a_19972_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3906 a_24092_5512# a_24004_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3907 vccd1 a_23833_25200# a_23728_25244# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X3908 a_21336_23589# a_5539_23589# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X3909 vccd1 a_11628_18056# a_13776_18100# vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3910 a_24540_11784# a_24452_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3911 vccd1 a_17820_18056# a_17732_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3912 vccd1 a_7190_18884# a_7646_19438# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3913 vccd1 a_13900_5079# a_13812_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3914 a_26780_3511# a_26692_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3915 vccd1 a_9408_25940# DIGITAL_OUT[0] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3916 vccd1 a_22972_22760# a_22884_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3917 a_14372_18884# a_4815_20408# a_14188_18884# vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3918 a_12856_16620# a_12455_16576# a_11799_16488# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3919 a_9176_16177# a_9076_15704# a_8972_16177# vccd1 pfet_06v0 ad=0.58035p pd=2.155u as=0.2847p ps=1.615u w=1.095u l=0.5u
X3920 a_26108_16488# a_26020_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3921 a_3619_17272# a_3949_17272# a_4069_17316# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3922 vccd1 a_8156_17584# a_6328_17342# vccd1 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3923 vssd1 a_19556_23992# a_20260_23588# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3924 vccd1 a_10676_16152# a_11919_14964# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3925 vssd1 a_4569_12176# a_4464_12316# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3926 a_19164_19624# a_19076_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3927 vccd1 a_20956_7080# a_20868_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3928 a_5732_22804# a_5612_23118# vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X3929 vssd1 a_6271_22596# a_6747_22020# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3930 a_27116_19191# a_27028_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3931 a_13984_13884# a_11872_13467# a_13672_13884# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3932 vccd1 a_2052_25940# a_9408_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3933 a_4233_23152# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X3934 a_27116_16055# a_27028_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3935 a_17820_3944# a_17732_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3936 a_2444_24328# a_7259_24800# vccd1 vccd1 pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
X3937 a_14986_14964# a_9532_13685# a_14092_14920# vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3938 a_9900_13396# a_9444_13880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X3939 SDAC[6] a_1772_23544# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3940 a_4731_20872# a_5019_20408# a_4935_20452# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X3941 a_3207_19288# a_3479_18840# a_3228_17317# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3942 a_13452_5079# a_13364_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3943 a_20508_8648# a_20420_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3944 vccd1 a_6383_25940# a_6839_25962# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3945 vssd1 a_6383_21028# a_6859_20452# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3946 a_27452_7080# a_27364_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3947 a_17680_23676# a_15568_23992# a_17368_23676# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3948 SDAC[5] a_1772_20408# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3949 a_23084_8215# a_22996_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3950 a_4233_18448# a_3816_18588# a_4609_18588# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3951 vccd1 a_12543_14964# a_12999_14986# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3952 a_1772_9432# a_3564_9432# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3953 vssd1 a_23725_24904# a_23845_24948# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3954 vccd1 a_11884_5079# a_11796_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3955 a_1772_6296# a_3564_6296# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3956 vccd1 a_4573_11000# a_4693_11620# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3957 a_5237_19669# a_4233_20016# vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3958 a_14012_3944# a_13924_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3959 a_1772_3160# a_3564_3160# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3960 a_13538_11828# a_12854_11828# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X3961 a_8004_24856# a_7884_24328# vssd1 vssd1 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3962 vssd1 a_5836_22760# a_10820_20452# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X3963 vccd1 a_21292_9783# a_21204_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3964 a_26220_6647# a_26132_6744# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3965 vccd1 a_21292_6647# a_21204_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3966 vccd1 a_2140_17302# a_7281_7142# vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3967 a_14538_13016# a_2140_17302# a_14350_13016# vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3968 vssd1 a_3564_20408# a_1772_20408# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D129 vssd1 a_3072_10564# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3969 DIGITAL_OUT[2] a_17024_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3970 a_8009_22804# a_7279_22826# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X3971 a_12984_21324# a_12432_21307# a_12780_21324# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3972 a_11961_25200# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X3973 vssd1 a_7055_22804# a_7531_23379# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3974 vccd1 a_15804_3944# a_15716_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3975 a_26108_22327# a_26020_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3976 a_23196_19624# a_23108_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3977 a_11628_18056# a_13496_17337# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3978 vssd1 a_9900_24756# a_9812_24856# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3979 a_9699_17396# a_9559_17540# a_9211_17272# vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X3980 a_10876_5512# a_10788_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3981 vssd1 a_24640_25940# DIGITAL_OUT[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3982 a_13780_18884# a_4815_20408# a_13604_18884# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X3983 a_2772_15052# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X3984 vssd1 a_6239_12568# a_6175_12613# vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3985 DIGITAL_OUT[1] a_13216_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3986 vccd1 a_3564_23544# a_1772_23544# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3987 a_6060_5079# a_5972_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3988 a_7134_10836# a_6470_10260# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3989 a_16192_25244# a_14576_25200# a_15064_25502# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3990 a_13496_17337# CLK vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3991 a_19052_11351# a_18964_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3992 vccd1 a_3564_20408# a_1772_20408# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3993 a_8568_7930# a_8752_8648# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.151p ps=1.185u w=0.36u l=0.6u
X3994 a_5627_23544# a_5975_23812# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X3995 vccd1 a_24540_3511# a_24452_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3996 a_5986_19460# a_5530_18884# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3997 vccd1 a_16588_8215# a_16500_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3998 vccd1 a_22188_19191# a_22100_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3999 vssd1 a_8568_7930# a_3564_6296# vssd1 nfet_06v0 ad=0.151p pd=1.185u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4000 a_20196_25940# a_19748_26471# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X4001 a_25212_19624# a_25124_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4002 vccd1 a_19164_16488# a_19076_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4003 vccd1 a_17859_24373# a_19748_26471# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X4004 a_2164_21236# a_1716_21767# vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X4005 a_15568_23992# a_15156_23671# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4006 a_23084_20759# a_22996_20856# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4007 vccd1 a_5836_22760# a_9444_19668# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4008 vccd1 a_20060_8648# a_19972_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4009 a_26556_16488# a_26468_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4010 vccd1 a_20060_5512# a_19972_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4011 a_17785_23632# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X4012 vccd1 a_20508_19624# a_20420_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4013 a_11936_17404# a_10320_17360# a_10808_17662# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4014 a_10808_13880# a_10136_13396# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X4015 vccd1 a_8412_3944# a_8324_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4016 a_6098_10260# a_5642_10260# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4017 a_27564_19191# a_27476_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4018 a_9360_11132# a_7744_11088# a_8232_11390# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4019 a_6215_25940# a_5759_25940# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4020 vccd1 a_2052_25940# a_9408_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4021 vccd1 a_4481_24757# a_11451_16488# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X4022 vssd1 a_26243_24765# a_22604_21976# vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4023 a_20299_21720# a_8009_22804# a_6060_23118# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4024 a_27564_16055# a_27476_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4025 vccd1 a_26556_8648# a_26468_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4026 vssd1 a_3542_22242# a_3682_22020# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4027 a_16364_16055# a_16276_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4028 vccd1 a_26556_5512# a_26468_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4029 a_17932_5079# a_17844_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4030 vccd1 a_27228_3511# a_27140_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4031 a_3484_5512# a_3396_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4032 a_10452_18840# a_16744_22042# vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X4033 vssd1 a_13496_15774# a_11548_13824# vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4034 a_23084_14487# a_22996_14584# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D130 a_1692_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4035 a_27564_8215# a_27476_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4036 a_4965_14136# a_1996_11000# a_5844_9880# vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4037 a_18716_8648# a_18628_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4038 a_23084_11351# a_22996_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4039 vccd1 a_1692_26427# a_8671_22020# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4040 a_14348_9783# a_14260_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4041 vccd1 a_3072_10564# a_12412_10348# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4042 vccd1 a_24004_22804# a_24640_25940# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4043 a_10428_7080# a_10340_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4044 vccd1 a_4815_20408# a_14736_20156# vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4045 vccd1 a_5948_3511# a_5860_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4046 DIGITAL_OUT[1] a_13216_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4047 vccd1 a_25212_22760# a_25124_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4048 vccd1 a_7259_24800# a_9444_19668# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4049 vccd1 a_23196_16488# a_23108_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4050 vccd1 a_15356_7080# a_15268_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4051 vccd1 a_25772_9783# a_25684_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4052 a_13292_21280# a_12984_21324# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4053 a_5767_12613# a_4964_9880# vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4054 vccd1 a_22636_17623# a_22548_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4055 vccd1 a_25772_6647# a_25684_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4056 a_11324_19624# a_11348_22065# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X4057 vccd1 a_3564_9432# a_1772_9432# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4058 vssd1 a_3072_10564# a_3024_18588# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4059 vccd1 a_3564_6296# a_1772_6296# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4060 DIGITAL_OUT[0] a_9408_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4061 a_6060_23118# a_8009_22804# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4062 a_11248_20452# a_5836_22760# vssd1 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4063 vccd1 a_10472_14181# a_5724_9432# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4064 vccd1 a_3564_3160# a_1772_3160# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4065 a_26556_22327# a_26468_22424# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4066 vccd1 a_20060_19191# a_19972_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4067 vccd1 a_18403_23197# a_13820_23544# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4068 vccd1 a_25212_16488# a_25124_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4069 a_22748_3944# a_22660_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4070 a_9479_10261# a_8121_13016# a_7820_7564# vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4071 vccd1 a_3816_18588# a_4233_18448# vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X4072 a_13496_17337# CLK vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4073 a_20396_16055# a_20308_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4074 a_13608_19712# a_13120_20112# a_13868_19756# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4075 vccd1 a_11772_3944# a_11684_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4076 a_13452_8648# a_13364_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4077 a_21404_16488# a_21316_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4078 a_25660_19624# a_25572_19668# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4079 a_3036_7080# a_2948_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4080 a_5577_9040# a_5160_9180# a_5953_9180# vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X4081 vssd1 a_4731_20872# a_17499_24856# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4082 vccd1 a_24540_8648# a_24452_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4083 DIGITAL_OUT[2] a_17024_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4084 vccd1 a_24540_5512# a_24452_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4085 a_15632_25244# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X4086 vccd1 a_6388_6390# a_2220_24686# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4087 a_18847_24460# a_17947_24328# vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X4088 SDAC[6] a_1772_23544# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4089 vccd1 a_20956_19624# a_20868_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4090 a_10903_10216# a_11664_10704# a_11455_10348# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X4091 vssd1 a_10732_24328# a_10684_24856# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X4092 a_7337_20856# a_6607_20452# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X4093 vccd1 a_15244_10216# a_15156_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4094 a_12104_20452# a_5836_22760# vssd1 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4095 a_6531_15357# a_6861_15429# a_6981_15539# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X4096 a_12732_13440# a_12424_13484# vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X4097 vccd1 a_9211_17272# a_9123_17317# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4098 vccd1 a_6553_24373# a_6431_22804# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4099 a_12108_21664# a_15456_19368# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X4100 vccd1 a_1916_17302# a_8736_19363# vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
D131 a_3072_10564# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4101 a_10871_12268# a_13910_11850# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X4102 vssd1 a_4481_24757# a_6115_23668# vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X4103 vccd1 a_13496_17337# a_11628_18056# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4104 a_17820_16488# a_17732_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4105 vccd1 a_24428_20759# a_24340_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4106 vccd1 a_4380_3944# a_4292_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4107 a_18828_9783# a_18740_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4108 vccd1 a_24640_25940# DIGITAL_OUT[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D132 a_5940_6390# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4109 a_14908_7080# a_14820_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4110 SDAC[2] a_1772_9432# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4111 vccd1 a_10540_5079# a_10452_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4112 SDAC[1] a_1772_6296# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4113 DIGITAL_OUT[1] a_13216_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4114 DIGITAL_OUT[4] a_21392_25940# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4115 vssd1 a_25648_25560# EOC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4116 vccd1 a_25660_22760# a_25572_22804# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4117 a_19648_21976# a_6553_24373# vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X4118 a_15848_20128# a_5237_19669# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X4119 a_14092_14920# a_9532_13685# vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X4120 vssd1 a_3564_9432# a_1772_9432# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4121 vccd1 a_7055_22804# a_7511_22826# vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4122 vssd1 a_1916_22021# a_1828_22065# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4123 SDAC[0] a_1772_3160# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4124 a_20956_8648# a_20868_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4125 a_13815_25380# a_14471_25571# a_14367_25615# vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4126 a_9127_22596# a_8671_22020# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4127 vccd1 a_11961_12656# a_11856_12700# vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4128 a_6154_19460# a_5530_18884# a_5986_19460# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
D133 a_1692_17302# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4129 vssd1 a_19357_18632# a_19477_18676# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4130 vccd1 a_12189_14136# a_12309_14756# vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4131 DIGITAL_OUT[0] a_9408_25940# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4132 a_9559_17540# a_10320_17360# a_10111_17775# vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X4133 a_18716_13352# a_18628_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4134 a_18403_18493# a_18733_18565# a_18853_18675# vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X4135 vccd1 a_24428_14487# a_24340_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4136 a_6844_3511# a_6756_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4137 a_14460_3944# a_14372_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4138 a_18716_10216# a_18628_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4139 vccd1 a_24428_11351# a_24340_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4140 a_23833_25200# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X4141 vccd1 a_25660_16488# a_25572_16532# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4142 a_10092_5079# a_10004_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4143 a_2876_22848# a_2568_22892# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4144 a_24092_7080# a_24004_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4145 vssd1 a_3072_10564# a_7952_9564# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4146 vccd1 a_7068_3944# a_6980_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4147 a_8225_19669# a_2164_21236# a_7932_20453# vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4148 a_7605_15540# a_7485_15496# a_6861_15429# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X4149 a_2016_13467# a_1604_13880# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4150 a_10808_13396# a_9076_15704# a_10808_13880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4151 a_6266_10260# a_5642_10260# a_6098_10260# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4152 a_2016_10331# a_1604_10744# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4153 vccd1 a_2444_24328# a_2340_24372# vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4154 vccd1 a_27004_13352# a_26916_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4155 a_20060_11784# a_19972_11828# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4156 a_2568_18188# a_1604_18584# a_2364_18188# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4157 a_21852_16488# a_21764_16532# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4158 a_26668_12919# a_26580_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4159 a_16588_5079# a_16500_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4160 vccd1 a_15244_8215# a_15156_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4161 a_4116_8780# a_2948_9176# a_3912_8780# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4162 vccd1 a_21516_18056# a_21428_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4163 vccd1 a_18256_25560# DIGITAL_OUT[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4164 vccd1 a_2444_26249# COMP_CLK vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4165 a_9744_8392# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4166 a_2876_13440# a_2568_13484# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4167 a_21628_21192# a_21540_21236# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4168 vssd1 a_4573_14136# a_4693_14180# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4169 a_2876_10304# a_2568_10348# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4170 a_9744_13016# a_9332_12695# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4171 vccd1 a_9644_5079# a_9556_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4172 vccd1 a_6266_10260# a_6702_10260# vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4173 a_15916_11351# a_15828_11448# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4174 vssd1 a_4573_11000# a_4693_11044# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4175 a_22748_13352# a_22660_13396# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4176 vccd1 a_15692_10216# a_15604_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4177 vssd1 a_17024_25940# DIGITAL_OUT[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4178 a_3524_24460# a_3404_24812# vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4179 vssd1 a_11548_13824# a_11460_13880# vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X4180 a_22748_10216# a_22660_10260# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4181 a_11043_10748# a_10903_10216# a_10555_10216# vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X4182 a_8225_19669# a_3703_18840# vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4183 a_21740_17623# a_21652_17720# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4184 vccd1 a_25212_8648# a_25124_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4185 a_17605_20452# a_2052_19288# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4186 vccd1 a_17820_7080# a_17732_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4187 a_1692_8215# a_1604_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4188 SDAC[2] a_1772_9432# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4189 a_2444_26249# a_4236_26254# vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4190 vssd1 a_8132_24372# a_8836_24372# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4191 vccd1 a_17632_21976# a_5019_20408# vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4192 vccd1 a_25212_5512# a_25124_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4193 vccd1 a_21180_3511# a_21092_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4194 a_2140_5512# a_2052_5556# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4195 a_4836_19288# a_4716_18840# a_2220_14136# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4196 a_19164_14920# a_19076_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4197 vccd1 a_19724_12919# a_19636_13016# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4198 a_14908_3511# a_14820_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4199 vccd1 a_24876_20759# a_24788_20856# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4200 vccd1 a_13496_17337# a_11628_18056# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4201 vccd1 a_8860_3944# a_8772_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4202 a_9196_5079# a_9108_5176# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4203 a_26220_8215# a_26132_8312# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4204 vccd1 a_4604_6647# a_4516_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4205 vssd1 a_25648_25560# EOC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4206 vssd1 a_6172_9432# a_5636_9476# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4207 a_13518_12404# a_12854_11828# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4208 vccd1 a_13496_15774# a_11548_13824# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4209 vccd1 a_4604_3511# a_4516_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4210 vccd1 a_27676_3511# a_27588_3608# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4211 a_2772_15052# a_1604_15448# a_2568_15052# vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4212 vccd1 a_3932_5512# a_3844_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4213 vccd1 a_14012_7080# a_13924_7124# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4214 vssd1 a_3004_21664# a_2940_21720# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4215 a_7485_13928# a_5573_11829# vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4216 vccd1 a_1692_18528# a_9332_25239# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4217 a_2772_19756# a_3072_10564# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X4218 a_10876_7080# a_10788_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4219 a_14796_9783# a_14708_9880# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4220 vssd1 a_4716_25204# a_4628_25248# vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4221 a_7792_23676# a_4481_24757# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X4222 a_13831_22596# a_13375_22020# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4223 a_19052_16055# a_18964_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4224 vccd1 a_24876_14487# a_24788_14584# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4225 vccd1 a_4380_5079# a_4292_5176# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4226 vssd1 a_6563_11784# a_6431_11828# vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X4227 vccd1 a_23196_8648# a_23108_8692# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4228 a_7042_19460# a_6358_19378# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X4229 vccd1 a_23196_5512# a_23108_5556# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4230 vccd1 a_24876_11351# a_24788_11448# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4231 a_12533_10052# a_12413_9432# a_11789_9432# vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4232 vccd1 a_21336_23589# a_4236_26254# vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4233 vssd1 a_3564_15704# a_1772_15704# vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D134 vssd1 a_4481_24757# diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4234 a_25212_24328# a_25124_24372# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4235 a_2940_21720# a_2820_21192# a_2672_21782# vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X4236 a_21404_3944# a_21316_3988# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4237 vssd1 a_8232_11390# a_8040_11503# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X4238 vccd1 a_18268_19191# a_18180_19288# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4239 a_23196_14920# a_23108_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4240 vccd1 a_27452_13352# a_27364_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4241 a_6944_9880# a_6532_9559# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4242 vccd1 a_25324_17623# a_25236_17720# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4243 vccd1 a_27116_9783# a_27028_9880# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4244 a_2364_15052# a_2264_15008# vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4245 vccd1 a_19724_8215# a_19636_8312# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4246 a_11664_10704# a_11548_13824# vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4247 vccd1 a_27116_6647# a_27028_6744# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4248 vccd1 a_19612_19624# a_19524_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4249 vccd1 a_21964_18056# a_21876_18100# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4250 vccd1 a_1692_10688# a_9332_12695# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4251 DIGITAL_OUT[3] a_18256_25560# vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4252 a_16709_21720# a_14953_22424# vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4253 a_3004_21664# a_7259_24800# vccd1 vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4254 a_6383_21028# a_5759_20452# a_6215_21028# vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4255 a_11968_23292# a_9856_22875# a_11656_23292# vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X4256 a_25212_18056# a_25124_18100# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4257 vccd1 a_6328_17342# a_1692_10688# vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4258 a_25212_14920# a_25124_14964# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4259 a_8644_14181# a_4348_7909# vssd1 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4260 a_24004_22804# a_23556_23335# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X4261 a_23084_19191# a_22996_19288# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4262 a_3484_7080# a_3396_7124# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4263 vssd1 a_17024_25940# DIGITAL_OUT[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4264 a_3972_24860# a_3136_24443# a_3728_24460# vssd1 nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4265 a_23084_16055# a_22996_16152# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4266 a_17932_12919# a_17844_13016# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4267 vccd1 a_9920_20096# a_4815_20408# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4268 vccd1 a_13116_3944# a_13028_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4269 a_1692_10688# a_6328_17342# vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X4270 a_18312_22021# a_2276_22424# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X4271 a_4481_24757# a_10192_8692# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4272 a_15288_22021# a_12308_22020# vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X4273 vccd1 a_14649_21584# a_14544_21724# vccd1 pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4274 a_2856_13884# a_2016_13467# a_2568_13484# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4275 a_6495_21724# a_3072_10564# a_5895_21372# vssd1 nfet_06v0 ad=86.399994f pd=0.84u as=0.1989p ps=1.465u w=0.36u l=0.6u
X4276 a_5612_23118# a_14953_22424# vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4277 a_2856_10748# a_2016_10331# a_2568_10348# vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4278 vssd1 a_6060_23118# a_5524_23288# vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4279 a_8156_17584# a_9800_18056# vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4280 a_16588_8648# a_16500_8692# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4281 vssd1 a_1772_9432# SDAC[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4282 a_6235_20452# a_5759_20452# vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4283 vccd1 a_23644_19624# a_23556_19668# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4284 vssd1 a_8156_17584# a_6440_18056# vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4285 a_21653_23379# a_21533_23269# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X4286 vssd1 a_15064_12613# a_8300_8648# vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X4287 vccd1 a_1692_18528# a_1604_18584# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4288 a_2016_17720# a_1916_17302# a_1812_17720# vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4289 a_4069_17870# a_3949_17272# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4290 a_3324_16576# a_3016_16620# vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4291 vccd1 a_26108_10216# a_26020_10260# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4292 a_23221_24947# a_23101_24837# vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X4293 a_6935_21724# a_5895_21372# vssd1 vssd1 nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4294 vccd1 a_4481_24757# a_13868_19756# vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4295 vccd1 a_9532_3944# a_9444_3988# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D135 a_2220_24686# vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4296 vccd1 a_1692_10688# a_1604_15448# vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4297 a_4069_14734# a_3949_14136# vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4298 a_15392_13824# a_14652_12605# vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X4299 a_1792_16532# a_1692_16488# vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4300 a_13494_14136# a_8519_13836# vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X4301 a_5500_3511# a_5412_3608# vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4302 vccd1 a_14708_18100# a_15456_19368# vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X4303 vccd1 a_22300_13352# a_22212_13396# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4304 a_9540_12268# a_9532_13685# a_10180_11828# vccd1 pfet_06v0 ad=0.2464p pd=2u as=0.1736p ps=1.18u w=0.56u l=0.5u
X4305 vccd1 a_27116_23895# a_27028_23992# vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4306 vssd1 a_3072_10564# a_3472_17020# vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4307 a_12628_13484# a_4481_24757# vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
.ends

